-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    num_cont : in  std_logic_vector(15 downto 0);
    row1 : in  std_logic_vector(15 downto 0);
    col1 : in  std_logic_vector(15 downto 0);
    rk1 : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 96)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal num_cont_buffer :  std_logic_vector(15 downto 0);
  signal num_cont_update_enable: Boolean;
  signal row1_buffer :  std_logic_vector(15 downto 0);
  signal row1_update_enable: Boolean;
  signal col1_buffer :  std_logic_vector(15 downto 0);
  signal col1_update_enable: Boolean;
  signal rk1_buffer :  std_logic_vector(15 downto 0);
  signal rk1_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_45_branch_req_0 : boolean;
  signal phi_stmt_47_req_1 : boolean;
  signal phi_stmt_47_req_0 : boolean;
  signal phi_stmt_47_ack_0 : boolean;
  signal n_address_281_51_buf_req_0 : boolean;
  signal n_address_281_51_buf_ack_0 : boolean;
  signal n_address_281_51_buf_req_1 : boolean;
  signal n_address_281_51_buf_ack_1 : boolean;
  signal phi_stmt_52_req_1 : boolean;
  signal phi_stmt_52_req_0 : boolean;
  signal phi_stmt_52_ack_0 : boolean;
  signal n_word_start_270_57_buf_req_0 : boolean;
  signal n_word_start_270_57_buf_ack_0 : boolean;
  signal n_word_start_270_57_buf_req_1 : boolean;
  signal n_word_start_270_57_buf_ack_1 : boolean;
  signal n_winr_210_71_buf_req_0 : boolean;
  signal n_winr_210_71_buf_ack_0 : boolean;
  signal n_winr_210_71_buf_req_1 : boolean;
  signal phi_stmt_58_req_0 : boolean;
  signal phi_stmt_58_req_1 : boolean;
  signal phi_stmt_58_ack_0 : boolean;
  signal n_left_289_60_buf_req_0 : boolean;
  signal n_left_289_60_buf_ack_0 : boolean;
  signal n_left_289_60_buf_req_1 : boolean;
  signal n_left_289_60_buf_ack_1 : boolean;
  signal nl_start_36_61_buf_req_0 : boolean;
  signal nl_start_36_61_buf_ack_0 : boolean;
  signal nl_start_36_61_buf_req_1 : boolean;
  signal nl_start_36_61_buf_ack_1 : boolean;
  signal phi_stmt_62_req_0 : boolean;
  signal phi_stmt_62_req_1 : boolean;
  signal phi_stmt_62_ack_0 : boolean;
  signal n_blk_309_64_buf_req_0 : boolean;
  signal n_blk_309_64_buf_ack_0 : boolean;
  signal n_blk_309_64_buf_req_1 : boolean;
  signal n_blk_309_64_buf_ack_1 : boolean;
  signal type_cast_66_inst_req_0 : boolean;
  signal type_cast_66_inst_ack_0 : boolean;
  signal type_cast_66_inst_req_1 : boolean;
  signal type_cast_66_inst_ack_1 : boolean;
  signal phi_stmt_67_req_1 : boolean;
  signal phi_stmt_67_req_0 : boolean;
  signal phi_stmt_67_ack_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_req_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_ack_0 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_req_1 : boolean;
  signal W_c3_165_delayed_14_0_171_inst_ack_1 : boolean;
  signal n_winr_210_71_buf_ack_1 : boolean;
  signal phi_stmt_72_req_0 : boolean;
  signal phi_stmt_72_req_1 : boolean;
  signal phi_stmt_72_ack_0 : boolean;
  signal n_col_223_74_buf_req_0 : boolean;
  signal n_col_223_74_buf_ack_0 : boolean;
  signal n_col_223_74_buf_req_1 : boolean;
  signal n_col_223_74_buf_ack_1 : boolean;
  signal phi_stmt_77_req_1 : boolean;
  signal phi_stmt_77_req_0 : boolean;
  signal phi_stmt_77_ack_0 : boolean;
  signal n_row_235_81_buf_req_0 : boolean;
  signal n_row_235_81_buf_ack_0 : boolean;
  signal n_row_235_81_buf_req_1 : boolean;
  signal n_row_235_81_buf_ack_1 : boolean;
  signal array_obj_ref_134_index_offset_req_0 : boolean;
  signal array_obj_ref_134_index_offset_ack_0 : boolean;
  signal array_obj_ref_134_index_offset_req_1 : boolean;
  signal array_obj_ref_134_index_offset_ack_1 : boolean;
  signal addr_of_135_final_reg_req_0 : boolean;
  signal addr_of_135_final_reg_ack_0 : boolean;
  signal addr_of_135_final_reg_req_1 : boolean;
  signal addr_of_135_final_reg_ack_1 : boolean;
  signal ptr_deref_139_load_0_req_0 : boolean;
  signal ptr_deref_139_load_0_ack_0 : boolean;
  signal ptr_deref_139_load_0_req_1 : boolean;
  signal ptr_deref_139_load_0_ack_1 : boolean;
  signal slice_143_inst_req_0 : boolean;
  signal slice_143_inst_ack_0 : boolean;
  signal slice_143_inst_req_1 : boolean;
  signal slice_143_inst_ack_1 : boolean;
  signal slice_147_inst_req_0 : boolean;
  signal slice_147_inst_ack_0 : boolean;
  signal slice_147_inst_req_1 : boolean;
  signal slice_147_inst_ack_1 : boolean;
  signal slice_151_inst_req_0 : boolean;
  signal slice_151_inst_ack_0 : boolean;
  signal slice_151_inst_req_1 : boolean;
  signal slice_151_inst_ack_1 : boolean;
  signal slice_155_inst_req_0 : boolean;
  signal slice_155_inst_ack_0 : boolean;
  signal slice_155_inst_req_1 : boolean;
  signal slice_155_inst_ack_1 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_req_0 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_ack_0 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_req_1 : boolean;
  signal W_c1_157_delayed_14_0_157_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_161_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_161_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_161_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_161_inst_ack_1 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_req_0 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_ack_0 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_req_1 : boolean;
  signal W_c2_161_delayed_14_0_164_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_168_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_168_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_168_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_168_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_175_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_175_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_175_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_175_inst_ack_1 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_req_0 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_ack_0 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_req_1 : boolean;
  signal W_c4_169_delayed_14_0_178_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_182_inst_req_0 : boolean;
  signal WPIPE_input_pipe1_182_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_182_inst_req_1 : boolean;
  signal WPIPE_input_pipe1_182_inst_ack_1 : boolean;
  signal do_while_stmt_45_branch_ack_0 : boolean;
  signal do_while_stmt_45_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 96) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= num_cont;
  num_cont_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= row1;
  row1_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= col1;
  col1_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(63 downto 48) <= rk1;
  rk1_buffer <= in_buffer_data_out(63 downto 48);
  in_buffer_data_in(79 downto 64) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(79 downto 64);
  in_buffer_data_in(95 downto 80) <= ct;
  ct_buffer <= in_buffer_data_out(95 downto 80);
  in_buffer_data_in(tag_length + 95 downto 96) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 95 downto 96);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(207 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_27/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/branch_block_stmt_27__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44__exit__
      -- CP-element group 0: 	 branch_block_stmt_27/do_while_stmt_45__entry__
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44/$entry
      -- CP-element group 0: 	 branch_block_stmt_27/assign_stmt_33_to_assign_stmt_44/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	207 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_27/$exit
      -- CP-element group 1: 	 branch_block_stmt_27/branch_block_stmt_27__exit__
      -- CP-element group 1: 	 branch_block_stmt_27/do_while_stmt_45__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(207);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_27/do_while_stmt_45/$entry
      -- CP-element group 2: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	207 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_27/do_while_stmt_45/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	205 
    -- CP-element group 5: 	206 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/condition_done
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	204 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_27/do_while_stmt_45/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(204);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	135 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	59 
    -- CP-element group 7: 	78 
    -- CP-element group 7: 	99 
    -- CP-element group 7: 	118 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	137 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	61 
    -- CP-element group 8: 	80 
    -- CP-element group 8: 	101 
    -- CP-element group 8: 	120 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	131 
    -- CP-element group 9: 	132 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	149 
    -- CP-element group 9: 	203 
    -- CP-element group 9: 	150 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	72 
    -- CP-element group 9: 	73 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	94 
    -- CP-element group 9: 	112 
    -- CP-element group 9: 	113 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	14 
    -- CP-element group 10: 	203 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_45_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(14) & access_T_CP_0_elements(203);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	131 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	112 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	114 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= access_T_CP_0_elements(131) & access_T_CP_0_elements(15) & access_T_CP_0_elements(34) & access_T_CP_0_elements(53) & access_T_CP_0_elements(72) & access_T_CP_0_elements(93) & access_T_CP_0_elements(112) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	133 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	75 
    -- CP-element group 12: 	96 
    -- CP-element group 12: 	115 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	204 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	131 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	53 
    -- CP-element group 12: 	72 
    -- CP-element group 12: 	93 
    -- CP-element group 12: 	112 
    -- CP-element group 12:  members (8) 
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(133) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(56) & access_T_CP_0_elements(75) & access_T_CP_0_elements(96) & access_T_CP_0_elements(115);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	132 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	54 
    -- CP-element group 13: 	73 
    -- CP-element group 13: 	94 
    -- CP-element group 13: 	113 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	57 
    -- CP-element group 13: 	76 
    -- CP-element group 13: 	97 
    -- CP-element group 13: 	116 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(132) & access_T_CP_0_elements(16) & access_T_CP_0_elements(35) & access_T_CP_0_elements(54) & access_T_CP_0_elements(73) & access_T_CP_0_elements(94) & access_T_CP_0_elements(113);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	134 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	77 
    -- CP-element group 14: 	98 
    -- CP-element group 14: 	117 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= access_T_CP_0_elements(134) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(58) & access_T_CP_0_elements(77) & access_T_CP_0_elements(98) & access_T_CP_0_elements(117);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	151 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: 	151 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resized_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/req
      -- 
    req_387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_134_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_loopback_sample_req_ps
      -- 
    phi_stmt_47_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_47_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_47_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_entry_sample_req_ps
      -- 
    phi_stmt_47_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_47_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_47_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_47_phi_mux_ack_ps
      -- 
    phi_stmt_47_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_47_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_update_start_
      -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_update_completed__ps
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_50_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(27), ack => access_T_CP_0_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(30), ack => n_address_281_51_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_update_start_
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => n_address_281_51_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_281_51_buf_ack_0, ack => access_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_address_51_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address_281_51_buf_ack_1, ack => access_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	177 
    -- CP-element group 35: 	184 
    -- CP-element group 35: 	191 
    -- CP-element group 35: 	198 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(177) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	175 
    -- CP-element group 39: 	182 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	189 
    -- CP-element group 39: 	196 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_loopback_sample_req_ps
      -- 
    phi_stmt_52_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_52_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_52_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_entry_sample_req_ps
      -- 
    phi_stmt_52_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_52_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_52_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_52_phi_mux_ack_ps
      -- 
    phi_stmt_52_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_52_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_start__ps
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_start__ps
      -- CP-element group 46: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_start_
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_completed__ps
      -- 
    access_T_CP_0_elements(47) <= access_T_CP_0_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_56_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(46), ack => access_T_CP_0_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_start__ps
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/req
      -- 
    req_115_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_115_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(49), ack => n_word_start_270_57_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_start_
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/req
      -- 
    req_120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(50), ack => n_word_start_270_57_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Sample/ack
      -- 
    ack_116_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_270_57_buf_ack_0, ack => access_T_CP_0_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_word_start_57_Update/ack
      -- 
    ack_121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_word_start_270_57_buf_ack_1, ack => access_T_CP_0_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	12 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	11 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_start_
      -- 
    access_T_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	13 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_start_
      -- 
    access_T_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(58);
      gj_access_T_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	11 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_start__ps
      -- 
    access_T_CP_0_elements(55) <= access_T_CP_0_elements(11);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	13 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(13);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	7 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_trigger
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(7);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_sample_req
      -- CP-element group 60: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_loopback_sample_req_ps
      -- 
    phi_stmt_58_loopback_sample_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_58_loopback_sample_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(60), ack => phi_stmt_58_req_0); -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(8);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_sample_req
      -- CP-element group 62: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_entry_sample_req_ps
      -- 
    phi_stmt_58_entry_sample_req_135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_58_entry_sample_req_135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_58_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_phi_mux_ack
      -- CP-element group 63: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_58_phi_mux_ack_ps
      -- 
    phi_stmt_58_phi_mux_ack_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_58_ack_0, ack => access_T_CP_0_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_start__ps
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/req
      -- 
    req_151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => n_left_289_60_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_start__ps
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_start_
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/req
      -- 
    req_156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(65), ack => n_left_289_60_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Sample/ack
      -- 
    ack_152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_289_60_buf_ack_0, ack => access_T_CP_0_elements(66)); -- 
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_left_60_Update/ack
      -- 
    ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_left_289_60_buf_ack_1, ack => access_T_CP_0_elements(67)); -- 
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(68), ack => nl_start_36_61_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_start_
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(69), ack => nl_start_36_61_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_36_61_buf_ack_0, ack => access_T_CP_0_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_nl_start_61_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nl_start_36_61_buf_ack_1, ack => access_T_CP_0_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	9 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	12 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	11 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_start_
      -- 
    access_T_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	184 
    -- CP-element group 73: 	191 
    -- CP-element group 73: 	198 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	13 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_start_
      -- 
    access_T_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(184) & access_T_CP_0_elements(191) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	11 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_start__ps
      -- 
    access_T_CP_0_elements(74) <= access_T_CP_0_elements(11);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	12 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	13 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_start__ps
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(13);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	182 
    -- CP-element group 77: 	14 
    -- CP-element group 77: 	189 
    -- CP-element group 77: 	196 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	7 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_trigger
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(7);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_sample_req
      -- CP-element group 79: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_loopback_sample_req_ps
      -- 
    phi_stmt_62_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_62_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(79), ack => phi_stmt_62_req_0); -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	8 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_trigger
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(8);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_sample_req
      -- CP-element group 81: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_entry_sample_req_ps
      -- 
    phi_stmt_62_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_62_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => phi_stmt_62_req_1); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_phi_mux_ack
      -- CP-element group 82: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_62_phi_mux_ack_ps
      -- 
    phi_stmt_62_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_62_ack_0, ack => access_T_CP_0_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_start__ps
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/req
      -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => n_blk_309_64_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_start__ps
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_start_
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/req
      -- 
    req_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(84), ack => n_blk_309_64_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Sample/ack
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_309_64_buf_ack_0, ack => access_T_CP_0_elements(85)); -- 
    -- CP-element group 86:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_completed__ps
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_blk_64_Update/ack
      -- 
    ack_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_blk_309_64_buf_ack_1, ack => access_T_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/rr
      -- 
    rr_223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(89), ack => type_cast_66_inst_req_0); -- 
    access_T_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(87) & access_T_CP_0_elements(91);
      gj_access_T_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_start_
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/cr
      -- 
    cr_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(90), ack => type_cast_66_inst_req_1); -- 
    access_T_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(88) & access_T_CP_0_elements(92);
      gj_access_T_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (4) 
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_completed__ps
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Sample/ra
      -- 
    ra_224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_0, ack => access_T_CP_0_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_66_Update/ca
      -- 
    ca_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_66_inst_ack_1, ack => access_T_CP_0_elements(92)); -- 
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	11 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_start_
      -- 
    access_T_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	9 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	98 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	13 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_start_
      -- 
    access_T_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(98);
      gj_access_T_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(11);
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	12 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	13 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_start__ps
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(13);
    -- CP-element group 98:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	14 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	94 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	7 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(7);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_sample_req
      -- CP-element group 100: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_loopback_sample_req_ps
      -- 
    phi_stmt_67_loopback_sample_req_240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_loopback_sample_req_240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_67_req_1); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	8 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_trigger
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(8);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_sample_req
      -- CP-element group 102: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_entry_sample_req_ps
      -- 
    phi_stmt_67_entry_sample_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_67_entry_sample_req_243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => phi_stmt_67_req_0); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_phi_mux_ack
      -- CP-element group 103: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_67_phi_mux_ack_ps
      -- 
    phi_stmt_67_phi_mux_ack_246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_67_ack_0, ack => access_T_CP_0_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_start_
      -- 
    -- Element group access_T_CP_0_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	107 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_completed__ps
      -- 
    access_T_CP_0_elements(106) <= access_T_CP_0_elements(107);
    -- CP-element group 107:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	106 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_70_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(107) is a control-delay.
    cp_element_107_delay: control_delay_element  generic map(name => " 107_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(105), ack => access_T_CP_0_elements(107), clk => clk, reset =>reset);
    -- CP-element group 108:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/req
      -- CP-element group 108: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_start__ps
      -- 
    req_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(108), ack => n_winr_210_71_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_start_
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/req
      -- 
    req_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(109), ack => n_winr_210_71_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (4) 
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_completed__ps
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Sample/ack
      -- 
    ack_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_210_71_buf_ack_0, ack => access_T_CP_0_elements(110)); -- 
    -- CP-element group 111:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (4) 
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_completed__ps
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_winr_71_Update/ack
      -- 
    ack_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_winr_210_71_buf_ack_1, ack => access_T_CP_0_elements(111)); -- 
    -- CP-element group 112:  join  transition  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	9 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	12 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	11 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_start_
      -- 
    access_T_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	9 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	117 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	13 
    -- CP-element group 113:  members (1) 
      -- CP-element group 113: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_start_
      -- 
    access_T_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(117);
      gj_access_T_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	11 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_start__ps
      -- 
    access_T_CP_0_elements(114) <= access_T_CP_0_elements(11);
    -- CP-element group 115:  join  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	12 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(115) is bound as output of CP function.
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	13 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_start__ps
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(13);
    -- CP-element group 117:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	14 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	113 
    -- CP-element group 117:  members (2) 
      -- CP-element group 117: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_completed_
      -- CP-element group 117: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	7 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_trigger
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(7);
    -- CP-element group 119:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_sample_req
      -- CP-element group 119: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_loopback_sample_req_ps
      -- 
    phi_stmt_72_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(119), ack => phi_stmt_72_req_0); -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	8 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_trigger
      -- 
    access_T_CP_0_elements(120) <= access_T_CP_0_elements(8);
    -- CP-element group 121:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_sample_req
      -- CP-element group 121: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_entry_sample_req_ps
      -- 
    phi_stmt_72_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_72_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(121), ack => phi_stmt_72_req_1); -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (2) 
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_phi_mux_ack
      -- CP-element group 122: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_72_phi_mux_ack_ps
      -- 
    phi_stmt_72_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_72_ack_0, ack => access_T_CP_0_elements(122)); -- 
    -- CP-element group 123:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (4) 
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_start__ps
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/req
      -- 
    req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(123), ack => n_col_223_74_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (4) 
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_start__ps
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_start_
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(124), ack => n_col_223_74_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(124) is bound as output of CP function.
    -- CP-element group 125:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_completed__ps
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Sample/ack
      -- 
    ack_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_223_74_buf_ack_0, ack => access_T_CP_0_elements(125)); -- 
    -- CP-element group 126:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_completed__ps
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_col_74_Update/ack
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_223_74_buf_ack_1, ack => access_T_CP_0_elements(126)); -- 
    -- CP-element group 127:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_start__ps
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(127) is bound as output of CP function.
    -- CP-element group 128:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (2) 
      -- CP-element group 128: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_start__ps
      -- CP-element group 128: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_start_
      -- 
    -- Element group access_T_CP_0_elements(128) is bound as output of CP function.
    -- CP-element group 129:  join  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	130 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_completed__ps
      -- 
    access_T_CP_0_elements(129) <= access_T_CP_0_elements(130);
    -- CP-element group 130:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	129 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_76_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(130) is a control-delay.
    cp_element_130_delay: control_delay_element  generic map(name => " 130_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(128), ack => access_T_CP_0_elements(130), clk => clk, reset =>reset);
    -- CP-element group 131:  join  transition  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	9 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	12 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	11 
    -- CP-element group 131:  members (1) 
      -- CP-element group 131: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_start_
      -- 
    access_T_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	9 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	13 
    -- CP-element group 132:  members (1) 
      -- CP-element group 132: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_start_
      -- 
    access_T_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	12 
    -- CP-element group 133:  members (1) 
      -- CP-element group 133: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(133) is bound as output of CP function.
    -- CP-element group 134:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	14 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(134) is bound as output of CP function.
    -- CP-element group 135:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	7 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_trigger
      -- 
    access_T_CP_0_elements(135) <= access_T_CP_0_elements(7);
    -- CP-element group 136:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (2) 
      -- CP-element group 136: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_sample_req
      -- CP-element group 136: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_loopback_sample_req_ps
      -- 
    phi_stmt_77_loopback_sample_req_328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_77_loopback_sample_req_328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(136), ack => phi_stmt_77_req_1); -- 
    -- Element group access_T_CP_0_elements(136) is bound as output of CP function.
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	8 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_trigger
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(8);
    -- CP-element group 138:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138:  members (2) 
      -- CP-element group 138: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_sample_req
      -- CP-element group 138: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_entry_sample_req_ps
      -- 
    phi_stmt_77_entry_sample_req_331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_77_entry_sample_req_331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(138), ack => phi_stmt_77_req_0); -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (2) 
      -- CP-element group 139: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_phi_mux_ack
      -- CP-element group 139: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/phi_stmt_77_phi_mux_ack_ps
      -- 
    phi_stmt_77_phi_mux_ack_334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_77_ack_0, ack => access_T_CP_0_elements(139)); -- 
    -- CP-element group 140:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_sample_start__ps
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_sample_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_sample_start_
      -- CP-element group 140: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (2) 
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_update_start__ps
      -- CP-element group 141: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_update_start_
      -- 
    -- Element group access_T_CP_0_elements(141) is bound as output of CP function.
    -- CP-element group 142:  join  transition  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	143 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (1) 
      -- CP-element group 142: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_update_completed__ps
      -- 
    access_T_CP_0_elements(142) <= access_T_CP_0_elements(143);
    -- CP-element group 143:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/type_cast_80_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(143) is a control-delay.
    cp_element_143_delay: control_delay_element  generic map(name => " 143_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(141), ack => access_T_CP_0_elements(143), clk => clk, reset =>reset);
    -- CP-element group 144:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (4) 
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_sample_start__ps
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_sample_start_
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Sample/$entry
      -- CP-element group 144: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Sample/req
      -- 
    req_355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => n_row_235_81_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (4) 
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_update_start__ps
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_update_start_
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Update/$entry
      -- CP-element group 145: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Update/req
      -- 
    req_360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(145), ack => n_row_235_81_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(145) is bound as output of CP function.
    -- CP-element group 146:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Sample/ack
      -- 
    ack_356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_235_81_buf_ack_0, ack => access_T_CP_0_elements(146)); -- 
    -- CP-element group 147:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (4) 
      -- CP-element group 147: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_update_completed__ps
      -- CP-element group 147: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/R_n_row_81_Update/ack
      -- 
    ack_361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_235_81_buf_ack_1, ack => access_T_CP_0_elements(147)); -- 
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	152 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	153 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	153 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_sample_start_
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/$entry
      -- CP-element group 148: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/req
      -- 
    req_402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(148), ack => addr_of_135_final_reg_req_0); -- 
    access_T_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(152) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	9 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	157 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	154 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_update_start_
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/$entry
      -- CP-element group 149: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/req
      -- 
    req_407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(149), ack => addr_of_135_final_reg_req_1); -- 
    access_T_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	9 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_update_start
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/req
      -- 
    req_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => array_obj_ref_134_index_offset_req_1); -- 
    access_T_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(153);
      gj_access_T_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	20 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	204 
    -- CP-element group 151: marked-successors 
    -- CP-element group 151: 	16 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_sample_complete
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Sample/ack
      -- 
    ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_134_index_offset_ack_0, ack => access_T_CP_0_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	148 
    -- CP-element group 152:  members (8) 
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_root_address_calculated
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_offset_calculated
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_final_index_sum_regn_Update/ack
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/$entry
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/$exit
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/sum_rename_req
      -- CP-element group 152: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/array_obj_ref_134_base_plus_offset/sum_rename_ack
      -- 
    ack_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_134_index_offset_ack_1, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	148 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/$exit
      -- CP-element group 153: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_request/ack
      -- 
    ack_403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_135_final_reg_ack_0, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	149 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (19) 
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/addr_of_135_complete/ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_root_address_calculated
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_address_resized
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/base_resize_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_addr_resize/base_resize_ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/sum_rename_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_base_plus_offset/sum_rename_ack
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/$entry
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/$exit
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/root_register_req
      -- CP-element group 154: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_word_addrgen/root_register_ack
      -- 
    ack_408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_135_final_reg_ack_1, ack => access_T_CP_0_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (5) 
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/$entry
      -- CP-element group 155: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/rr
      -- 
    rr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(155), ack => ptr_deref_139_load_0_req_0); -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(154) & access_T_CP_0_elements(157);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	173 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	169 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (5) 
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_update_start_
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/$entry
      -- CP-element group 156: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/cr
      -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(156), ack => ptr_deref_139_load_0_req_1); -- 
    access_T_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(173) & access_T_CP_0_elements(161) & access_T_CP_0_elements(165) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	149 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (5) 
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/$exit
      -- CP-element group 157: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Sample/word_access_start/word_0/ra
      -- 
    ra_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_load_0_ack_0, ack => access_T_CP_0_elements(157)); -- 
    -- CP-element group 158:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	171 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	163 
    -- CP-element group 158: 	167 
    -- CP-element group 158:  members (9) 
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/word_access_complete/word_0/ca
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/$entry
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/$exit
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/merge_req
      -- CP-element group 158: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/ptr_deref_139_Update/ptr_deref_139_Merge/merge_ack
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_139_load_0_ack_1, ack => access_T_CP_0_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/rr
      -- 
    rr_466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(159), ack => slice_143_inst_req_0); -- 
    access_T_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(161);
      gj_access_T_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	180 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_update_start_
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/cr
      -- 
    cr_471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(160), ack => slice_143_inst_req_1); -- 
    access_T_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	156 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Sample/ra
      -- 
    ra_467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_143_inst_ack_0, ack => access_T_CP_0_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	179 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_143_Update/ca
      -- 
    ca_472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_143_inst_ack_1, ack => access_T_CP_0_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	158 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/rr
      -- 
    rr_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => slice_147_inst_req_0); -- 
    access_T_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(165);
      gj_access_T_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	187 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_update_start_
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/cr
      -- 
    cr_485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(164), ack => slice_147_inst_req_1); -- 
    access_T_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	156 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Sample/ra
      -- 
    ra_481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_0, ack => access_T_CP_0_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	186 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_147_Update/ca
      -- 
    ca_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_147_inst_ack_1, ack => access_T_CP_0_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	158 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/rr
      -- 
    rr_494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(167), ack => slice_151_inst_req_0); -- 
    access_T_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(169);
      gj_access_T_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	194 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_update_start_
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/cr
      -- 
    cr_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(168), ack => slice_151_inst_req_1); -- 
    access_T_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	156 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Sample/ra
      -- 
    ra_495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_0, ack => access_T_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	193 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_151_Update/ca
      -- 
    ca_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_151_inst_ack_1, ack => access_T_CP_0_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	158 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/rr
      -- 
    rr_508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(171), ack => slice_155_inst_req_0); -- 
    access_T_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(158) & access_T_CP_0_elements(173);
      gj_access_T_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	201 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_update_start_
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/cr
      -- 
    cr_513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(172), ack => slice_155_inst_req_1); -- 
    access_T_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	156 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Sample/ra
      -- 
    ra_509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_0, ack => access_T_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	200 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/$exit
      -- CP-element group 174: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/slice_155_Update/ca
      -- 
    ca_514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_155_inst_ack_1, ack => access_T_CP_0_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	39 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/req
      -- 
    req_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(175), ack => W_c1_157_delayed_14_0_157_inst_req_0); -- 
    access_T_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(177);
      gj_access_T_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	180 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_update_start_
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/req
      -- 
    req_527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(176), ack => W_c1_157_delayed_14_0_157_inst_req_1); -- 
    access_T_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(180);
      gj_access_T_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: 	35 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Sample/ack
      -- 
    ack_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_157_delayed_14_0_157_inst_ack_0, ack => access_T_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_159_Update/ack
      -- 
    ack_528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c1_157_delayed_14_0_157_inst_ack_1, ack => access_T_CP_0_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: 	162 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	202 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/req
      -- 
    req_536_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_536_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(179), ack => WPIPE_input_pipe1_161_inst_req_0); -- 
    access_T_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(178) & access_T_CP_0_elements(162) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	176 
    -- CP-element group 180: 	160 
    -- CP-element group 180:  members (6) 
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_update_start_
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Sample/ack
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/req
      -- 
    ack_537_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_161_inst_ack_0, ack => access_T_CP_0_elements(180)); -- 
    req_541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => WPIPE_input_pipe1_161_inst_req_1); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	186 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_161_Update/ack
      -- 
    ack_542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_161_inst_ack_1, ack => access_T_CP_0_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	39 
    -- CP-element group 182: 	77 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/req
      -- 
    req_550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => W_c2_161_delayed_14_0_164_inst_req_0); -- 
    access_T_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(77) & access_T_CP_0_elements(184);
      gj_access_T_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	187 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_update_start_
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/req
      -- 
    req_555_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_555_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(183), ack => W_c2_161_delayed_14_0_164_inst_req_1); -- 
    access_T_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(187);
      gj_access_T_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: 	35 
    -- CP-element group 184: 	73 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Sample/ack
      -- 
    ack_551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_161_delayed_14_0_164_inst_ack_0, ack => access_T_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_166_Update/ack
      -- 
    ack_556_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c2_161_delayed_14_0_164_inst_ack_1, ack => access_T_CP_0_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	181 
    -- CP-element group 186: 	185 
    -- CP-element group 186: 	166 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/req
      -- 
    req_564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(186), ack => WPIPE_input_pipe1_168_inst_req_0); -- 
    access_T_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(181) & access_T_CP_0_elements(185) & access_T_CP_0_elements(166) & access_T_CP_0_elements(188);
      gj_access_T_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	183 
    -- CP-element group 187: 	164 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_update_start_
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Sample/ack
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/req
      -- 
    ack_565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_168_inst_ack_0, ack => access_T_CP_0_elements(187)); -- 
    req_569_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_569_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(187), ack => WPIPE_input_pipe1_168_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	193 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_168_Update/ack
      -- 
    ack_570_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_168_inst_ack_1, ack => access_T_CP_0_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	39 
    -- CP-element group 189: 	77 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/req
      -- 
    req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(189), ack => W_c3_165_delayed_14_0_171_inst_req_0); -- 
    access_T_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(77) & access_T_CP_0_elements(191);
      gj_access_T_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_update_start_
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/req
      -- 
    req_583_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_583_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => W_c3_165_delayed_14_0_171_inst_req_1); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(194);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	35 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	73 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Sample/ack
      -- 
    ack_579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_165_delayed_14_0_171_inst_ack_0, ack => access_T_CP_0_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_173_Update/ack
      -- 
    ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c3_165_delayed_14_0_171_inst_ack_1, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	170 
    -- CP-element group 193: 	188 
    -- CP-element group 193: 	192 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/req
      -- 
    req_592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(193), ack => WPIPE_input_pipe1_175_inst_req_0); -- 
    access_T_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(170) & access_T_CP_0_elements(188) & access_T_CP_0_elements(192) & access_T_CP_0_elements(195);
      gj_access_T_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	168 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_update_start_
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/req
      -- 
    ack_593_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_175_inst_ack_0, ack => access_T_CP_0_elements(194)); -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(194), ack => WPIPE_input_pipe1_175_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	200 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_175_Update/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_175_inst_ack_1, ack => access_T_CP_0_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	39 
    -- CP-element group 196: 	77 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/req
      -- 
    req_606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(196), ack => W_c4_169_delayed_14_0_178_inst_req_0); -- 
    access_T_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(39) & access_T_CP_0_elements(77) & access_T_CP_0_elements(198);
      gj_access_T_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_update_start_
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/req
      -- 
    req_611_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_611_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(197), ack => W_c4_169_delayed_14_0_178_inst_req_1); -- 
    access_T_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(201);
      gj_access_T_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	35 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	73 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Sample/ack
      -- 
    ack_607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_169_delayed_14_0_178_inst_ack_0, ack => access_T_CP_0_elements(198)); -- 
    -- CP-element group 199:  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/assign_stmt_180_Update/ack
      -- 
    ack_612_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_c4_169_delayed_14_0_178_inst_ack_1, ack => access_T_CP_0_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	174 
    -- CP-element group 200: 	195 
    -- CP-element group 200: 	199 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/req
      -- 
    req_620_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_620_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(200), ack => WPIPE_input_pipe1_182_inst_req_0); -- 
    access_T_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= access_T_CP_0_elements(174) & access_T_CP_0_elements(195) & access_T_CP_0_elements(199) & access_T_CP_0_elements(202);
      gj_access_T_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	172 
    -- CP-element group 201: 	197 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_update_start_
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/req
      -- 
    ack_621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_182_inst_ack_0, ack => access_T_CP_0_elements(201)); -- 
    req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => WPIPE_input_pipe1_182_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	179 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/WPIPE_input_pipe1_182_Update/ack
      -- 
    ack_626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_182_inst_ack_1, ack => access_T_CP_0_elements(202)); -- 
    -- CP-element group 203:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	9 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	10 
    -- CP-element group 203:  members (1) 
      -- CP-element group 203: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(203) is a control-delay.
    cp_element_203_delay: control_delay_element  generic map(name => " 203_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(203), clk => clk, reset =>reset);
    -- CP-element group 204:  join  transition  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	12 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	151 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	6 
    -- CP-element group 204:  members (1) 
      -- CP-element group 204: 	 branch_block_stmt_27/do_while_stmt_45/do_while_stmt_45_loop_body/$exit
      -- 
    access_T_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(12) & access_T_CP_0_elements(202) & access_T_CP_0_elements(151);
      gj_access_T_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	5 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (2) 
      -- CP-element group 205: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/$exit
      -- CP-element group 205: 	 branch_block_stmt_27/do_while_stmt_45/loop_exit/ack
      -- 
    ack_631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_45_branch_ack_0, ack => access_T_CP_0_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	5 
    -- CP-element group 206: successors 
    -- CP-element group 206:  members (2) 
      -- CP-element group 206: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/$exit
      -- CP-element group 206: 	 branch_block_stmt_27/do_while_stmt_45/loop_taken/ack
      -- 
    ack_635_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_45_branch_ack_1, ack => access_T_CP_0_elements(206)); -- 
    -- CP-element group 207:  transition  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	3 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	1 
    -- CP-element group 207:  members (1) 
      -- CP-element group 207: 	 branch_block_stmt_27/do_while_stmt_45/$exit
      -- 
    access_T_CP_0_elements(207) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_45_terminator_636: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_45_terminator_636", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(206),loop_terminate => access_T_CP_0_elements(205),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_47_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(33);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_47_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_47_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_52_phi_seq_122_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(45);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(47);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(51);
      access_T_CP_0_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(52);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_52_phi_seq_122 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_52_phi_seq_122") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_58_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(59);
      access_T_CP_0_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(67);
      access_T_CP_0_elements(60) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(70);
      access_T_CP_0_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(71);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_58_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_58_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(55), 
          phi_sample_ack => access_T_CP_0_elements(56), 
          phi_update_req => access_T_CP_0_elements(57), 
          phi_update_ack => access_T_CP_0_elements(58), 
          phi_mux_ack => access_T_CP_0_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_62_phi_seq_230_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(78);
      access_T_CP_0_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(85);
      access_T_CP_0_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(86);
      access_T_CP_0_elements(79) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(80);
      access_T_CP_0_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(92);
      access_T_CP_0_elements(81) <= phi_mux_reqs(1);
      phi_stmt_62_phi_seq_230 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_62_phi_seq_230") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(74), 
          phi_sample_ack => access_T_CP_0_elements(75), 
          phi_update_req => access_T_CP_0_elements(76), 
          phi_update_ack => access_T_CP_0_elements(77), 
          phi_mux_ack => access_T_CP_0_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_67_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(101);
      access_T_CP_0_elements(104)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(104);
      access_T_CP_0_elements(105)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(102) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(108)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(110);
      access_T_CP_0_elements(109)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(111);
      access_T_CP_0_elements(100) <= phi_mux_reqs(1);
      phi_stmt_67_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_67_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(95), 
          phi_sample_ack => access_T_CP_0_elements(96), 
          phi_update_req => access_T_CP_0_elements(97), 
          phi_update_ack => access_T_CP_0_elements(98), 
          phi_mux_ack => access_T_CP_0_elements(103), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_72_phi_seq_318_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(118);
      access_T_CP_0_elements(123)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(125);
      access_T_CP_0_elements(124)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(126);
      access_T_CP_0_elements(119) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(120);
      access_T_CP_0_elements(127)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(128)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(129);
      access_T_CP_0_elements(121) <= phi_mux_reqs(1);
      phi_stmt_72_phi_seq_318 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_72_phi_seq_318") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(114), 
          phi_sample_ack => access_T_CP_0_elements(115), 
          phi_update_req => access_T_CP_0_elements(116), 
          phi_update_ack => access_T_CP_0_elements(117), 
          phi_mux_ack => access_T_CP_0_elements(122), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_77_phi_seq_362_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(137);
      access_T_CP_0_elements(140)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(140);
      access_T_CP_0_elements(141)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(142);
      access_T_CP_0_elements(138) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(135);
      access_T_CP_0_elements(144)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(145)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(147);
      access_T_CP_0_elements(136) <= phi_mux_reqs(1);
      phi_stmt_77_phi_seq_362 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_77_phi_seq_362") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(133), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(134), 
          phi_mux_ack => access_T_CP_0_elements(139), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_126_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_206_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_219_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_232_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_242_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_294_wire : std_logic_vector(15 downto 0);
    signal ADD_u64_u64_279_wire : std_logic_vector(63 downto 0);
    signal AND_u1_u1_108_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_115_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_214_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_228_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_229_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_95_wire : std_logic_vector(0 downto 0);
    signal AND_u32_u32_261_wire : std_logic_vector(31 downto 0);
    signal EQ_u2_u1_104_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_111_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_118_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_91_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_98_wire : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_275_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_241_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_243_wire : std_logic_vector(15 downto 0);
    signal MUL_u16_u16_31_wire : std_logic_vector(15 downto 0);
    signal MUL_u32_u32_250_wire : std_logic_vector(31 downto 0);
    signal MUX_207_wire : std_logic_vector(15 downto 0);
    signal MUX_220_wire : std_logic_vector(15 downto 0);
    signal MUX_301_wire : std_logic_vector(15 downto 0);
    signal MUX_307_wire : std_logic_vector(15 downto 0);
    signal NEQ_u16_u1_313_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_119_wire : std_logic_vector(0 downto 0);
    signal R_address_133_resized : std_logic_vector(13 downto 0);
    signal R_address_133_scaled : std_logic_vector(13 downto 0);
    signal SUB_u16_u16_287_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_299_wire : std_logic_vector(15 downto 0);
    signal UGT_u16_u1_107_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_114_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_296_wire : std_logic_vector(0 downto 0);
    signal UGT_u16_u1_94_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_304_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_40_wire : std_logic_vector(0 downto 0);
    signal address_47 : std_logic_vector(63 downto 0);
    signal array_obj_ref_134_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_134_root_address : std_logic_vector(13 downto 0);
    signal c1_157_delayed_14_0_159 : std_logic_vector(0 downto 0);
    signal c1_87 : std_logic_vector(0 downto 0);
    signal c2_100 : std_logic_vector(0 downto 0);
    signal c2_161_delayed_14_0_166 : std_logic_vector(0 downto 0);
    signal c3_121 : std_logic_vector(0 downto 0);
    signal c3_165_delayed_14_0_173 : std_logic_vector(0 downto 0);
    signal c4_129 : std_logic_vector(0 downto 0);
    signal c4_169_delayed_14_0_180 : std_logic_vector(0 downto 0);
    signal col_72 : std_logic_vector(15 downto 0);
    signal col_done_199 : std_logic_vector(0 downto 0);
    signal fetch_addr_136 : std_logic_vector(31 downto 0);
    signal flag1_189 : std_logic_vector(0 downto 0);
    signal fn_blk_44 : std_logic_vector(15 downto 0);
    signal konst_103_wire_constant : std_logic_vector(1 downto 0);
    signal konst_106_wire_constant : std_logic_vector(15 downto 0);
    signal konst_110_wire_constant : std_logic_vector(1 downto 0);
    signal konst_113_wire_constant : std_logic_vector(15 downto 0);
    signal konst_117_wire_constant : std_logic_vector(1 downto 0);
    signal konst_127_wire_constant : std_logic_vector(15 downto 0);
    signal konst_203_wire_constant : std_logic_vector(15 downto 0);
    signal konst_205_wire_constant : std_logic_vector(15 downto 0);
    signal konst_216_wire_constant : std_logic_vector(15 downto 0);
    signal konst_218_wire_constant : std_logic_vector(15 downto 0);
    signal konst_231_wire_constant : std_logic_vector(15 downto 0);
    signal konst_260_wire_constant : std_logic_vector(31 downto 0);
    signal konst_268_wire_constant : std_logic_vector(1 downto 0);
    signal konst_274_wire_constant : std_logic_vector(31 downto 0);
    signal konst_278_wire_constant : std_logic_vector(63 downto 0);
    signal konst_295_wire_constant : std_logic_vector(15 downto 0);
    signal konst_297_wire_constant : std_logic_vector(15 downto 0);
    signal konst_303_wire_constant : std_logic_vector(15 downto 0);
    signal konst_306_wire_constant : std_logic_vector(15 downto 0);
    signal konst_39_wire_constant : std_logic_vector(15 downto 0);
    signal konst_42_wire_constant : std_logic_vector(15 downto 0);
    signal konst_85_wire_constant : std_logic_vector(1 downto 0);
    signal konst_90_wire_constant : std_logic_vector(1 downto 0);
    signal konst_93_wire_constant : std_logic_vector(15 downto 0);
    signal konst_97_wire_constant : std_logic_vector(1 downto 0);
    signal m_factor_33 : std_logic_vector(31 downto 0);
    signal n_address_281 : std_logic_vector(63 downto 0);
    signal n_address_281_51_buffered : std_logic_vector(63 downto 0);
    signal n_blk_309 : std_logic_vector(15 downto 0);
    signal n_blk_309_64_buffered : std_logic_vector(15 downto 0);
    signal n_col_223 : std_logic_vector(15 downto 0);
    signal n_col_223_74_buffered : std_logic_vector(15 downto 0);
    signal n_left_289 : std_logic_vector(15 downto 0);
    signal n_left_289_60_buffered : std_logic_vector(15 downto 0);
    signal n_row_235 : std_logic_vector(15 downto 0);
    signal n_row_235_81_buffered : std_logic_vector(15 downto 0);
    signal n_winr_210 : std_logic_vector(15 downto 0);
    signal n_winr_210_71_buffered : std_logic_vector(15 downto 0);
    signal n_word_start_270 : std_logic_vector(1 downto 0);
    signal n_word_start_270_57_buffered : std_logic_vector(1 downto 0);
    signal na1_245 : std_logic_vector(31 downto 0);
    signal na2_252 : std_logic_vector(31 downto 0);
    signal na3_257 : std_logic_vector(31 downto 0);
    signal na4_263 : std_logic_vector(15 downto 0);
    signal nl_start_36 : std_logic_vector(15 downto 0);
    signal nl_start_36_61_buffered : std_logic_vector(15 downto 0);
    signal num_blk_62 : std_logic_vector(15 downto 0);
    signal num_left_58 : std_logic_vector(15 downto 0);
    signal ptr_deref_139_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_139_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_139_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_139_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_139_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_77 : std_logic_vector(15 downto 0);
    signal type_cast_125_wire : std_logic_vector(15 downto 0);
    signal type_cast_249_wire : std_logic_vector(31 downto 0);
    signal type_cast_267_wire : std_logic_vector(1 downto 0);
    signal type_cast_276_wire : std_logic_vector(63 downto 0);
    signal type_cast_50_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_56_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_66_wire : std_logic_vector(15 downto 0);
    signal type_cast_70_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_76_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_80_wire_constant : std_logic_vector(15 downto 0);
    signal w1_144 : std_logic_vector(15 downto 0);
    signal w2_148 : std_logic_vector(15 downto 0);
    signal w3_152 : std_logic_vector(15 downto 0);
    signal w4_156 : std_logic_vector(15 downto 0);
    signal winr_67 : std_logic_vector(15 downto 0);
    signal winr_done_194 : std_logic_vector(0 downto 0);
    signal word_read_140 : std_logic_vector(63 downto 0);
    signal word_start_52 : std_logic_vector(1 downto 0);
    -- 
  begin -- 
    array_obj_ref_134_constant_part_of_offset <= "00000000000000";
    array_obj_ref_134_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_134_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_134_resized_base_address <= "00000000000000";
    konst_103_wire_constant <= "00";
    konst_106_wire_constant <= "0000000000000010";
    konst_110_wire_constant <= "01";
    konst_113_wire_constant <= "0000000000000001";
    konst_117_wire_constant <= "10";
    konst_127_wire_constant <= "0000000000000011";
    konst_203_wire_constant <= "0000000000000000";
    konst_205_wire_constant <= "0000000000000001";
    konst_216_wire_constant <= "0000000000000000";
    konst_218_wire_constant <= "0000000000000001";
    konst_231_wire_constant <= "0000000000000001";
    konst_260_wire_constant <= "00000000000000000000000000000011";
    konst_268_wire_constant <= "00";
    konst_274_wire_constant <= "00000000000000000000000000000010";
    konst_278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_295_wire_constant <= "0000000000000100";
    konst_297_wire_constant <= "0000000000000100";
    konst_303_wire_constant <= "0000000000000100";
    konst_306_wire_constant <= "0000000000000100";
    konst_39_wire_constant <= "0000000000000100";
    konst_42_wire_constant <= "0000000000000100";
    konst_85_wire_constant <= "00";
    konst_90_wire_constant <= "00";
    konst_93_wire_constant <= "0000000000000001";
    konst_97_wire_constant <= "01";
    ptr_deref_139_word_offset_0 <= "00000000000000";
    type_cast_50_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_56_wire_constant <= "00";
    type_cast_70_wire_constant <= "0000000000000000";
    type_cast_76_wire_constant <= "0000000000000000";
    type_cast_80_wire_constant <= "0000000000000000";
    phi_stmt_47: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_50_wire_constant & n_address_281_51_buffered;
      req <= phi_stmt_47_req_0 & phi_stmt_47_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_47",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_47_ack_0,
          idata => idata,
          odata => address_47,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_47
    phi_stmt_52: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_56_wire_constant & n_word_start_270_57_buffered;
      req <= phi_stmt_52_req_0 & phi_stmt_52_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_52",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_52_ack_0,
          idata => idata,
          odata => word_start_52,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_52
    phi_stmt_58: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_left_289_60_buffered & nl_start_36_61_buffered;
      req <= phi_stmt_58_req_0 & phi_stmt_58_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_58",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_58_ack_0,
          idata => idata,
          odata => num_left_58,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_58
    phi_stmt_62: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_blk_309_64_buffered & type_cast_66_wire;
      req <= phi_stmt_62_req_0 & phi_stmt_62_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_62",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_62_ack_0,
          idata => idata,
          odata => num_blk_62,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_62
    phi_stmt_67: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_70_wire_constant & n_winr_210_71_buffered;
      req <= phi_stmt_67_req_0 & phi_stmt_67_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_67",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_67_ack_0,
          idata => idata,
          odata => winr_67,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_67
    phi_stmt_72: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_col_223_74_buffered & type_cast_76_wire_constant;
      req <= phi_stmt_72_req_0 & phi_stmt_72_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_72",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_72_ack_0,
          idata => idata,
          odata => col_72,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_72
    phi_stmt_77: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_80_wire_constant & n_row_235_81_buffered;
      req <= phi_stmt_77_req_0 & phi_stmt_77_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_77",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_77_ack_0,
          idata => idata,
          odata => row_77,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_77
    -- flow-through select operator MUX_207_inst
    MUX_207_wire <= konst_203_wire_constant when (winr_done_194(0) /=  '0') else ADD_u16_u16_206_wire;
    -- flow-through select operator MUX_209_inst
    n_winr_210 <= MUX_207_wire when (flag1_189(0) /=  '0') else winr_67;
    -- flow-through select operator MUX_220_inst
    MUX_220_wire <= konst_216_wire_constant when (col_done_199(0) /=  '0') else ADD_u16_u16_219_wire;
    -- flow-through select operator MUX_222_inst
    n_col_223 <= MUX_220_wire when (AND_u1_u1_214_wire(0) /=  '0') else col_72;
    -- flow-through select operator MUX_234_inst
    n_row_235 <= ADD_u16_u16_232_wire when (AND_u1_u1_229_wire(0) /=  '0') else row_77;
    -- flow-through select operator MUX_269_inst
    n_word_start_270 <= type_cast_267_wire when (flag1_189(0) /=  '0') else konst_268_wire_constant;
    -- flow-through select operator MUX_280_inst
    n_address_281 <= type_cast_276_wire when (flag1_189(0) /=  '0') else ADD_u64_u64_279_wire;
    -- flow-through select operator MUX_288_inst
    n_left_289 <= nl_start_36 when (flag1_189(0) /=  '0') else SUB_u16_u16_287_wire;
    -- flow-through select operator MUX_301_inst
    MUX_301_wire <= SUB_u16_u16_299_wire when (UGT_u16_u1_296_wire(0) /=  '0') else fn_blk_44;
    -- flow-through select operator MUX_307_inst
    MUX_307_wire <= n_left_289 when (ULT_u16_u1_304_wire(0) /=  '0') else konst_306_wire_constant;
    -- flow-through select operator MUX_308_inst
    n_blk_309 <= MUX_301_wire when (flag1_189(0) /=  '0') else MUX_307_wire;
    -- flow-through select operator MUX_43_inst
    fn_blk_44 <= num_cont_buffer when (ULT_u16_u1_40_wire(0) /=  '0') else konst_42_wire_constant;
    slice_143_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_143_inst_req_0;
      slice_143_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_143_inst_req_1;
      slice_143_inst_ack_1<= update_ack(0);
      slice_143_inst: SliceSplitProtocol generic map(name => "slice_143_inst", in_data_width => 64, high_index => 63, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w1_144, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_147_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_147_inst_req_0;
      slice_147_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_147_inst_req_1;
      slice_147_inst_ack_1<= update_ack(0);
      slice_147_inst: SliceSplitProtocol generic map(name => "slice_147_inst", in_data_width => 64, high_index => 47, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w2_148, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_151_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_151_inst_req_0;
      slice_151_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_151_inst_req_1;
      slice_151_inst_ack_1<= update_ack(0);
      slice_151_inst: SliceSplitProtocol generic map(name => "slice_151_inst", in_data_width => 64, high_index => 31, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w3_152, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_155_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_155_inst_req_0;
      slice_155_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_155_inst_req_1;
      slice_155_inst_ack_1<= update_ack(0);
      slice_155_inst: SliceSplitProtocol generic map(name => "slice_155_inst", in_data_width => 64, high_index => 15, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => word_read_140, dout => w4_156, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_c1_157_delayed_14_0_157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c1_157_delayed_14_0_157_inst_req_0;
      W_c1_157_delayed_14_0_157_inst_ack_0<= wack(0);
      rreq(0) <= W_c1_157_delayed_14_0_157_inst_req_1;
      W_c1_157_delayed_14_0_157_inst_ack_1<= rack(0);
      W_c1_157_delayed_14_0_157_inst : InterlockBuffer generic map ( -- 
        name => "W_c1_157_delayed_14_0_157_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c1_87,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c1_157_delayed_14_0_159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c2_161_delayed_14_0_164_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c2_161_delayed_14_0_164_inst_req_0;
      W_c2_161_delayed_14_0_164_inst_ack_0<= wack(0);
      rreq(0) <= W_c2_161_delayed_14_0_164_inst_req_1;
      W_c2_161_delayed_14_0_164_inst_ack_1<= rack(0);
      W_c2_161_delayed_14_0_164_inst : InterlockBuffer generic map ( -- 
        name => "W_c2_161_delayed_14_0_164_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c2_100,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c2_161_delayed_14_0_166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c3_165_delayed_14_0_171_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c3_165_delayed_14_0_171_inst_req_0;
      W_c3_165_delayed_14_0_171_inst_ack_0<= wack(0);
      rreq(0) <= W_c3_165_delayed_14_0_171_inst_req_1;
      W_c3_165_delayed_14_0_171_inst_ack_1<= rack(0);
      W_c3_165_delayed_14_0_171_inst : InterlockBuffer generic map ( -- 
        name => "W_c3_165_delayed_14_0_171_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c3_121,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c3_165_delayed_14_0_173,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_c4_169_delayed_14_0_178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_c4_169_delayed_14_0_178_inst_req_0;
      W_c4_169_delayed_14_0_178_inst_ack_0<= wack(0);
      rreq(0) <= W_c4_169_delayed_14_0_178_inst_req_1;
      W_c4_169_delayed_14_0_178_inst_ack_1<= rack(0);
      W_c4_169_delayed_14_0_178_inst : InterlockBuffer generic map ( -- 
        name => "W_c4_169_delayed_14_0_178_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => c4_129,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => c4_169_delayed_14_0_180,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_nl_start_34_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := num_cont_buffer(15 downto 0);
      nl_start_36 <= tmp_var; -- 
    end process;
    addr_of_135_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_135_final_reg_req_0;
      addr_of_135_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_135_final_reg_req_1;
      addr_of_135_final_reg_ack_1<= rack(0);
      addr_of_135_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_135_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_134_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address_281_51_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address_281_51_buf_req_0;
      n_address_281_51_buf_ack_0<= wack(0);
      rreq(0) <= n_address_281_51_buf_req_1;
      n_address_281_51_buf_ack_1<= rack(0);
      n_address_281_51_buf : InterlockBuffer generic map ( -- 
        name => "n_address_281_51_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address_281,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address_281_51_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_blk_309_64_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_blk_309_64_buf_req_0;
      n_blk_309_64_buf_ack_0<= wack(0);
      rreq(0) <= n_blk_309_64_buf_req_1;
      n_blk_309_64_buf_ack_1<= rack(0);
      n_blk_309_64_buf : InterlockBuffer generic map ( -- 
        name => "n_blk_309_64_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_blk_309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_blk_309_64_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_223_74_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_223_74_buf_req_0;
      n_col_223_74_buf_ack_0<= wack(0);
      rreq(0) <= n_col_223_74_buf_req_1;
      n_col_223_74_buf_ack_1<= rack(0);
      n_col_223_74_buf : InterlockBuffer generic map ( -- 
        name => "n_col_223_74_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_223_74_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_left_289_60_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_left_289_60_buf_req_0;
      n_left_289_60_buf_ack_0<= wack(0);
      rreq(0) <= n_left_289_60_buf_req_1;
      n_left_289_60_buf_ack_1<= rack(0);
      n_left_289_60_buf : InterlockBuffer generic map ( -- 
        name => "n_left_289_60_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_left_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_left_289_60_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_235_81_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_235_81_buf_req_0;
      n_row_235_81_buf_ack_0<= wack(0);
      rreq(0) <= n_row_235_81_buf_req_1;
      n_row_235_81_buf_ack_1<= rack(0);
      n_row_235_81_buf : InterlockBuffer generic map ( -- 
        name => "n_row_235_81_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_235_81_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_winr_210_71_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_winr_210_71_buf_req_0;
      n_winr_210_71_buf_ack_0<= wack(0);
      rreq(0) <= n_winr_210_71_buf_req_1;
      n_winr_210_71_buf_ack_1<= rack(0);
      n_winr_210_71_buf : InterlockBuffer generic map ( -- 
        name => "n_winr_210_71_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_winr_210,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_winr_210_71_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_word_start_270_57_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_word_start_270_57_buf_req_0;
      n_word_start_270_57_buf_ack_0<= wack(0);
      rreq(0) <= n_word_start_270_57_buf_req_1;
      n_word_start_270_57_buf_ack_1<= rack(0);
      n_word_start_270_57_buf : InterlockBuffer generic map ( -- 
        name => "n_word_start_270_57_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_word_start_270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_word_start_270_57_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nl_start_36_61_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nl_start_36_61_buf_req_0;
      nl_start_36_61_buf_ack_0<= wack(0);
      rreq(0) <= nl_start_36_61_buf_req_1;
      nl_start_36_61_buf_ack_1<= rack(0);
      nl_start_36_61_buf : InterlockBuffer generic map ( -- 
        name => "nl_start_36_61_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nl_start_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nl_start_36_61_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_125_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := word_start_52(1 downto 0);
      type_cast_125_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_244_inst
    process(MUL_u16_u16_243_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_243_wire(15 downto 0);
      na1_245 <= tmp_var; -- 
    end process;
    -- interlock type_cast_249_inst
    process(n_winr_210) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_winr_210(15 downto 0);
      type_cast_249_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_251_inst
    process(MUL_u32_u32_250_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := MUL_u32_u32_250_wire(31 downto 0);
      na2_252 <= tmp_var; -- 
    end process;
    -- interlock type_cast_262_inst
    process(AND_u32_u32_261_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := AND_u32_u32_261_wire(15 downto 0);
      na4_263 <= tmp_var; -- 
    end process;
    -- interlock type_cast_267_inst
    process(na4_263) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 1 downto 0) := na4_263(1 downto 0);
      type_cast_267_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_276_inst
    process(LSHR_u32_u32_275_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_275_wire(31 downto 0);
      type_cast_276_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_32_inst
    process(MUL_u16_u16_31_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_31_wire(15 downto 0);
      m_factor_33 <= tmp_var; -- 
    end process;
    type_cast_66_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_66_inst_req_0;
      type_cast_66_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_66_inst_req_1;
      type_cast_66_inst_ack_1<= rack(0);
      type_cast_66_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_66_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_blk_44,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_66_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_134_index_1_rename
    process(R_address_133_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_address_133_resized;
      ov(13 downto 0) := iv;
      R_address_133_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_134_index_1_resize
    process(address_47) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := address_47;
      ov := iv(13 downto 0);
      R_address_133_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_134_root_address_inst
    process(array_obj_ref_134_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_134_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_134_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_addr_0
    process(ptr_deref_139_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_139_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_base_resize
    process(fetch_addr_136) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_136;
      ov := iv(13 downto 0);
      ptr_deref_139_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_gather_scatter
    process(ptr_deref_139_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_data_0;
      ov(63 downto 0) := iv;
      word_read_140 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_139_root_address_inst
    process(ptr_deref_139_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_139_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_139_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_45_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NEQ_u16_u1_313_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_45_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_45_branch_req_0,
          ack0 => do_while_stmt_45_branch_ack_0,
          ack1 => do_while_stmt_45_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_126_inst
    process(num_blk_62, type_cast_125_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_blk_62, type_cast_125_wire, tmp_var);
      ADD_u16_u16_126_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_206_inst
    process(winr_67) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(winr_67, konst_205_wire_constant, tmp_var);
      ADD_u16_u16_206_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_219_inst
    process(col_72) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_72, konst_218_wire_constant, tmp_var);
      ADD_u16_u16_219_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_232_inst
    process(row_77) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_77, konst_231_wire_constant, tmp_var);
      ADD_u16_u16_232_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_242_inst
    process(n_col_223, MUL_u16_u16_241_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(n_col_223, MUL_u16_u16_241_wire, tmp_var);
      ADD_u16_u16_242_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_294_inst
    process(fn_blk_44, na4_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(fn_blk_44, na4_263, tmp_var);
      ADD_u16_u16_294_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_256_inst
    process(na1_245, na2_252) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(na1_245, na2_252, tmp_var);
      na3_257 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_279_inst
    process(address_47) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address_47, konst_278_wire_constant, tmp_var);
      ADD_u64_u64_279_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_108_inst
    process(EQ_u2_u1_104_wire, UGT_u16_u1_107_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_104_wire, UGT_u16_u1_107_wire, tmp_var);
      AND_u1_u1_108_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_115_inst
    process(EQ_u2_u1_111_wire, UGT_u16_u1_114_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_111_wire, UGT_u16_u1_114_wire, tmp_var);
      AND_u1_u1_115_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_214_inst
    process(winr_done_194, flag1_189) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_194, flag1_189, tmp_var);
      AND_u1_u1_214_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_228_inst
    process(col_done_199, flag1_189) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_199, flag1_189, tmp_var);
      AND_u1_u1_228_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_229_inst
    process(winr_done_194, AND_u1_u1_228_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(winr_done_194, AND_u1_u1_228_wire, tmp_var);
      AND_u1_u1_229_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_95_inst
    process(EQ_u2_u1_91_wire, UGT_u16_u1_94_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_91_wire, UGT_u16_u1_94_wire, tmp_var);
      AND_u1_u1_95_wire <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_261_inst
    process(na3_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(na3_257, konst_260_wire_constant, tmp_var);
      AND_u32_u32_261_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_188_inst
    process(num_left_58, num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_left_58, num_blk_62, tmp_var);
      flag1_189 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_193_inst
    process(winr_67, rk1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(winr_67, rk1_buffer, tmp_var);
      winr_done_194 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_198_inst
    process(col_72, col1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_72, col1_buffer, tmp_var);
      col_done_199 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_104_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_103_wire_constant, tmp_var);
      EQ_u2_u1_104_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_111_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_110_wire_constant, tmp_var);
      EQ_u2_u1_111_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_118_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_117_wire_constant, tmp_var);
      EQ_u2_u1_118_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_86_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_85_wire_constant, tmp_var);
      c1_87 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_91_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_90_wire_constant, tmp_var);
      EQ_u2_u1_91_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_98_inst
    process(word_start_52) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(word_start_52, konst_97_wire_constant, tmp_var);
      EQ_u2_u1_98_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_275_inst
    process(na3_257) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(na3_257, konst_274_wire_constant, tmp_var);
      LSHR_u32_u32_275_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_241_inst
    process(ct_buffer, n_row_235) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, n_row_235, tmp_var);
      MUL_u16_u16_241_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_243_inst
    process(chl_in_buffer, ADD_u16_u16_242_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_in_buffer, ADD_u16_u16_242_wire, tmp_var);
      MUL_u16_u16_243_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_31_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_31_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_250_inst
    process(m_factor_33, type_cast_249_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(m_factor_33, type_cast_249_wire, tmp_var);
      MUL_u32_u32_250_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u16_u1_313_inst
    process(n_row_235, row1_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(n_row_235, row1_buffer, tmp_var);
      NEQ_u16_u1_313_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_119_inst
    process(AND_u1_u1_115_wire, EQ_u2_u1_118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_115_wire, EQ_u2_u1_118_wire, tmp_var);
      OR_u1_u1_119_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_120_inst
    process(AND_u1_u1_108_wire, OR_u1_u1_119_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_108_wire, OR_u1_u1_119_wire, tmp_var);
      c3_121 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_99_inst
    process(AND_u1_u1_95_wire, EQ_u2_u1_98_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_95_wire, EQ_u2_u1_98_wire, tmp_var);
      c2_100 <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_287_inst
    process(num_left_58, num_blk_62) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(num_left_58, num_blk_62, tmp_var);
      SUB_u16_u16_287_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u16_u16_299_inst
    process(konst_297_wire_constant, na4_263) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_297_wire_constant, na4_263, tmp_var);
      SUB_u16_u16_299_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_107_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_106_wire_constant, tmp_var);
      UGT_u16_u1_107_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_114_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_113_wire_constant, tmp_var);
      UGT_u16_u1_114_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_128_inst
    process(ADD_u16_u16_126_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_126_wire, konst_127_wire_constant, tmp_var);
      c4_129 <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_296_inst
    process(ADD_u16_u16_294_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ADD_u16_u16_294_wire, konst_295_wire_constant, tmp_var);
      UGT_u16_u1_296_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u16_u1_94_inst
    process(num_blk_62) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_blk_62, konst_93_wire_constant, tmp_var);
      UGT_u16_u1_94_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_304_inst
    process(n_left_289) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_left_289, konst_303_wire_constant, tmp_var);
      ULT_u16_u1_304_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_40_inst
    process(num_cont_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(num_cont_buffer, konst_39_wire_constant, tmp_var);
      ULT_u16_u1_40_wire <= tmp_var; --
    end process;
    -- shared split operator group (42) : array_obj_ref_134_index_offset 
    ApIntAdd_group_42: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_address_133_scaled;
      array_obj_ref_134_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_134_index_offset_req_0;
      array_obj_ref_134_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_134_index_offset_req_1;
      array_obj_ref_134_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_42_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_42_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_42",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared load operator group (0) : ptr_deref_139_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_139_load_0_req_0;
      ptr_deref_139_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_139_load_0_req_1;
      ptr_deref_139_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_139_word_address_0;
      ptr_deref_139_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_175_inst WPIPE_input_pipe1_168_inst WPIPE_input_pipe1_161_inst WPIPE_input_pipe1_182_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 3 downto 0);
      signal update_req, update_ack : BooleanArray( 3 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 3 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => true, 1 => true, 2 => true, 3 => true);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      sample_req_unguarded(3) <= WPIPE_input_pipe1_175_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_input_pipe1_168_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_input_pipe1_161_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_input_pipe1_182_inst_req_0;
      WPIPE_input_pipe1_175_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_input_pipe1_168_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_input_pipe1_161_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_input_pipe1_182_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(3) <= WPIPE_input_pipe1_175_inst_req_1;
      update_req_unguarded(2) <= WPIPE_input_pipe1_168_inst_req_1;
      update_req_unguarded(1) <= WPIPE_input_pipe1_161_inst_req_1;
      update_req_unguarded(0) <= WPIPE_input_pipe1_182_inst_req_1;
      WPIPE_input_pipe1_175_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_input_pipe1_168_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_input_pipe1_161_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_input_pipe1_182_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= c4_169_delayed_14_0_180(0);
      guard_vector(1)  <= c1_157_delayed_14_0_159(0);
      guard_vector(2)  <= c2_161_delayed_14_0_166(0);
      guard_vector(3)  <= c3_165_delayed_14_0_173(0);
      data_in <= w3_152 & w2_148 & w1_144 & w4_156;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 16, num_reqs => 4, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(95 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_1115_start: Boolean;
  signal convolution3D_CP_1115_symbol: Boolean;
  -- volatile/operator module components. 
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_649_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1339_inst_ack_1 : boolean;
  signal type_cast_665_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_req_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal type_cast_586_inst_req_1 : boolean;
  signal type_cast_573_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_0 : boolean;
  signal type_cast_645_inst_ack_0 : boolean;
  signal type_cast_598_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_ack_1 : boolean;
  signal type_cast_611_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_1 : boolean;
  signal type_cast_611_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_ack_0 : boolean;
  signal type_cast_623_inst_req_1 : boolean;
  signal type_cast_645_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_594_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_req_0 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal type_cast_623_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_ack_1 : boolean;
  signal type_cast_586_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_ack_1 : boolean;
  signal type_cast_548_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_ack_0 : boolean;
  signal type_cast_623_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_req_1 : boolean;
  signal type_cast_598_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_ack_1 : boolean;
  signal type_cast_623_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_569_inst_req_1 : boolean;
  signal type_cast_511_inst_req_0 : boolean;
  signal type_cast_523_inst_req_0 : boolean;
  signal type_cast_573_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_557_inst_req_0 : boolean;
  signal type_cast_665_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_ack_1 : boolean;
  signal type_cast_548_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_req_1 : boolean;
  signal type_cast_586_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_ack_1 : boolean;
  signal type_cast_665_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_619_inst_ack_0 : boolean;
  signal type_cast_511_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_req_0 : boolean;
  signal type_cast_665_inst_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal type_cast_598_inst_req_0 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_532_inst_req_0 : boolean;
  signal type_cast_1307_inst_ack_1 : boolean;
  signal if_stmt_673_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1303_inst_req_1 : boolean;
  signal type_cast_645_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_544_inst_ack_0 : boolean;
  signal type_cast_636_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_607_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_507_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_0 : boolean;
  signal type_cast_611_inst_req_1 : boolean;
  signal type_cast_536_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_582_inst_ack_1 : boolean;
  signal type_cast_598_inst_ack_0 : boolean;
  signal type_cast_511_inst_req_1 : boolean;
  signal type_cast_536_inst_ack_0 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_611_inst_ack_1 : boolean;
  signal type_cast_511_inst_ack_1 : boolean;
  signal type_cast_645_inst_req_1 : boolean;
  signal type_cast_1325_inst_ack_0 : boolean;
  signal type_cast_718_inst_req_0 : boolean;
  signal type_cast_1343_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_req_1 : boolean;
  signal type_cast_693_inst_req_1 : boolean;
  signal type_cast_1253_inst_ack_1 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal type_cast_548_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1339_inst_req_1 : boolean;
  signal type_cast_718_inst_ack_0 : boolean;
  signal type_cast_693_inst_req_0 : boolean;
  signal type_cast_693_inst_ack_0 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1303_inst_ack_0 : boolean;
  signal type_cast_693_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1236_inst_req_1 : boolean;
  signal type_cast_709_inst_req_0 : boolean;
  signal type_cast_709_inst_ack_0 : boolean;
  signal type_cast_548_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_1 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal if_stmt_673_branch_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_ack_1 : boolean;
  signal type_cast_709_inst_req_1 : boolean;
  signal type_cast_709_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_519_inst_req_0 : boolean;
  signal if_stmt_673_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1303_inst_req_0 : boolean;
  signal type_cast_586_inst_req_0 : boolean;
  signal addr_of_1233_final_reg_ack_1 : boolean;
  signal type_cast_1253_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_1 : boolean;
  signal type_cast_718_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1285_inst_ack_1 : boolean;
  signal type_cast_718_inst_ack_1 : boolean;
  signal type_cast_523_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1236_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_req_0 : boolean;
  signal type_cast_536_inst_ack_1 : boolean;
  signal type_cast_536_inst_req_1 : boolean;
  signal type_cast_523_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_ack_0 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_632_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1236_inst_req_0 : boolean;
  signal type_cast_523_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1267_inst_ack_0 : boolean;
  signal array_obj_ref_1232_index_offset_req_0 : boolean;
  signal type_cast_1325_inst_req_1 : boolean;
  signal type_cast_1289_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_444_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_444_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1236_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_444_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_444_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1303_inst_ack_1 : boolean;
  signal type_cast_1289_inst_ack_0 : boolean;
  signal type_cast_448_inst_req_0 : boolean;
  signal type_cast_448_inst_ack_0 : boolean;
  signal type_cast_1325_inst_ack_1 : boolean;
  signal type_cast_448_inst_req_1 : boolean;
  signal type_cast_448_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_457_inst_ack_1 : boolean;
  signal array_obj_ref_1232_index_offset_ack_0 : boolean;
  signal type_cast_461_inst_req_0 : boolean;
  signal type_cast_461_inst_ack_0 : boolean;
  signal type_cast_461_inst_req_1 : boolean;
  signal type_cast_461_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_469_inst_ack_1 : boolean;
  signal type_cast_473_inst_req_0 : boolean;
  signal type_cast_473_inst_ack_0 : boolean;
  signal type_cast_473_inst_req_1 : boolean;
  signal type_cast_473_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_482_inst_ack_1 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_494_inst_ack_1 : boolean;
  signal type_cast_498_inst_req_0 : boolean;
  signal type_cast_498_inst_ack_0 : boolean;
  signal type_cast_498_inst_req_1 : boolean;
  signal type_cast_498_inst_ack_1 : boolean;
  signal type_cast_1253_inst_ack_0 : boolean;
  signal type_cast_1325_inst_req_0 : boolean;
  signal type_cast_728_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1285_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_0 : boolean;
  signal type_cast_728_inst_req_1 : boolean;
  signal type_cast_728_inst_ack_1 : boolean;
  signal addr_of_1233_final_reg_req_1 : boolean;
  signal type_cast_1307_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1339_inst_ack_0 : boolean;
  signal type_cast_1253_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_ack_1 : boolean;
  signal array_obj_ref_763_index_offset_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1285_inst_ack_0 : boolean;
  signal array_obj_ref_763_index_offset_ack_0 : boolean;
  signal array_obj_ref_763_index_offset_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1285_inst_req_0 : boolean;
  signal array_obj_ref_763_index_offset_ack_1 : boolean;
  signal type_cast_1343_inst_req_1 : boolean;
  signal type_cast_1343_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_req_1 : boolean;
  signal addr_of_1233_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1339_inst_req_0 : boolean;
  signal addr_of_764_final_reg_req_0 : boolean;
  signal addr_of_764_final_reg_ack_0 : boolean;
  signal addr_of_764_final_reg_req_1 : boolean;
  signal addr_of_764_final_reg_ack_1 : boolean;
  signal addr_of_1233_final_reg_req_0 : boolean;
  signal type_cast_1307_inst_ack_0 : boolean;
  signal type_cast_1307_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_767_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_767_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_767_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_767_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1249_inst_req_0 : boolean;
  signal type_cast_771_inst_req_0 : boolean;
  signal type_cast_1271_inst_ack_1 : boolean;
  signal type_cast_771_inst_ack_0 : boolean;
  signal type_cast_771_inst_req_1 : boolean;
  signal type_cast_1271_inst_req_1 : boolean;
  signal type_cast_771_inst_ack_1 : boolean;
  signal type_cast_1289_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_780_inst_ack_1 : boolean;
  signal type_cast_1240_inst_ack_1 : boolean;
  signal type_cast_1240_inst_req_1 : boolean;
  signal type_cast_784_inst_req_0 : boolean;
  signal type_cast_1271_inst_ack_0 : boolean;
  signal type_cast_784_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_ack_1 : boolean;
  signal type_cast_784_inst_req_1 : boolean;
  signal type_cast_1271_inst_req_0 : boolean;
  signal type_cast_784_inst_ack_1 : boolean;
  signal type_cast_1289_inst_req_1 : boolean;
  signal array_obj_ref_1232_index_offset_ack_1 : boolean;
  signal type_cast_1343_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_798_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_798_inst_ack_0 : boolean;
  signal array_obj_ref_1232_index_offset_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_798_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_798_inst_ack_1 : boolean;
  signal type_cast_1240_inst_ack_0 : boolean;
  signal type_cast_1240_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1321_inst_req_1 : boolean;
  signal type_cast_802_inst_req_0 : boolean;
  signal type_cast_802_inst_ack_0 : boolean;
  signal type_cast_802_inst_req_1 : boolean;
  signal type_cast_802_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_816_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_816_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_816_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_816_inst_ack_1 : boolean;
  signal type_cast_754_inst_ack_0 : boolean;
  signal type_cast_1748_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1792_inst_req_1 : boolean;
  signal phi_stmt_986_ack_0 : boolean;
  signal type_cast_1758_inst_ack_1 : boolean;
  signal type_cast_820_inst_req_0 : boolean;
  signal type_cast_820_inst_ack_0 : boolean;
  signal type_cast_820_inst_req_1 : boolean;
  signal type_cast_820_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_834_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_834_inst_ack_0 : boolean;
  signal type_cast_1778_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_834_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1792_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_834_inst_ack_1 : boolean;
  signal type_cast_1778_inst_ack_0 : boolean;
  signal type_cast_838_inst_req_0 : boolean;
  signal type_cast_838_inst_ack_0 : boolean;
  signal type_cast_838_inst_req_1 : boolean;
  signal type_cast_838_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_852_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_852_inst_ack_0 : boolean;
  signal type_cast_1778_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_852_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_852_inst_ack_1 : boolean;
  signal type_cast_1778_inst_ack_1 : boolean;
  signal phi_stmt_993_ack_0 : boolean;
  signal type_cast_856_inst_req_0 : boolean;
  signal type_cast_856_inst_ack_0 : boolean;
  signal type_cast_856_inst_req_1 : boolean;
  signal type_cast_856_inst_ack_1 : boolean;
  signal type_cast_754_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_870_inst_req_0 : boolean;
  signal type_cast_754_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_870_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_870_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_870_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1795_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1795_inst_ack_0 : boolean;
  signal type_cast_874_inst_req_0 : boolean;
  signal type_cast_874_inst_ack_0 : boolean;
  signal type_cast_992_inst_req_0 : boolean;
  signal type_cast_874_inst_req_1 : boolean;
  signal type_cast_874_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_888_inst_ack_1 : boolean;
  signal type_cast_892_inst_req_0 : boolean;
  signal type_cast_892_inst_ack_0 : boolean;
  signal type_cast_1748_inst_req_1 : boolean;
  signal type_cast_892_inst_req_1 : boolean;
  signal phi_stmt_751_req_0 : boolean;
  signal type_cast_892_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1780_inst_req_0 : boolean;
  signal type_cast_1748_inst_ack_1 : boolean;
  signal ptr_deref_900_store_0_req_0 : boolean;
  signal ptr_deref_900_store_0_ack_0 : boolean;
  signal ptr_deref_900_store_0_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1795_inst_req_1 : boolean;
  signal ptr_deref_900_store_0_ack_1 : boolean;
  signal type_cast_948_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1795_inst_ack_1 : boolean;
  signal type_cast_948_inst_ack_0 : boolean;
  signal if_stmt_914_branch_req_0 : boolean;
  signal if_stmt_914_branch_ack_1 : boolean;
  signal if_stmt_914_branch_ack_0 : boolean;
  signal type_cast_992_inst_ack_0 : boolean;
  signal if_stmt_965_branch_req_0 : boolean;
  signal if_stmt_965_branch_ack_1 : boolean;
  signal if_stmt_965_branch_ack_0 : boolean;
  signal phi_stmt_751_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1014_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1014_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1014_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1014_inst_ack_1 : boolean;
  signal type_cast_1758_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1780_inst_ack_0 : boolean;
  signal type_cast_992_inst_req_1 : boolean;
  signal type_cast_1018_inst_req_0 : boolean;
  signal type_cast_1018_inst_ack_0 : boolean;
  signal type_cast_992_inst_ack_1 : boolean;
  signal type_cast_1018_inst_req_1 : boolean;
  signal type_cast_1018_inst_ack_1 : boolean;
  signal phi_stmt_986_req_1 : boolean;
  signal type_cast_1033_inst_req_0 : boolean;
  signal type_cast_1033_inst_ack_0 : boolean;
  signal type_cast_1033_inst_req_1 : boolean;
  signal type_cast_1033_inst_ack_1 : boolean;
  signal type_cast_1758_inst_ack_0 : boolean;
  signal if_stmt_1040_branch_req_0 : boolean;
  signal if_stmt_1040_branch_ack_1 : boolean;
  signal if_stmt_1040_branch_ack_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_0 : boolean;
  signal array_obj_ref_1079_index_offset_ack_0 : boolean;
  signal array_obj_ref_1079_index_offset_req_1 : boolean;
  signal array_obj_ref_1079_index_offset_ack_1 : boolean;
  signal addr_of_1080_final_reg_req_0 : boolean;
  signal addr_of_1080_final_reg_ack_0 : boolean;
  signal addr_of_1080_final_reg_req_1 : boolean;
  signal addr_of_1080_final_reg_ack_1 : boolean;
  signal ptr_deref_1083_store_0_req_0 : boolean;
  signal ptr_deref_1083_store_0_ack_0 : boolean;
  signal ptr_deref_1083_store_0_req_1 : boolean;
  signal ptr_deref_1083_store_0_ack_1 : boolean;
  signal type_cast_1090_inst_req_0 : boolean;
  signal type_cast_1090_inst_ack_0 : boolean;
  signal type_cast_1090_inst_req_1 : boolean;
  signal type_cast_1090_inst_ack_1 : boolean;
  signal type_cast_1094_inst_req_0 : boolean;
  signal type_cast_1094_inst_ack_0 : boolean;
  signal type_cast_1094_inst_req_1 : boolean;
  signal type_cast_1094_inst_ack_1 : boolean;
  signal type_cast_1098_inst_req_0 : boolean;
  signal type_cast_1098_inst_ack_0 : boolean;
  signal type_cast_1098_inst_req_1 : boolean;
  signal type_cast_1098_inst_ack_1 : boolean;
  signal type_cast_1102_inst_req_0 : boolean;
  signal type_cast_1102_inst_ack_0 : boolean;
  signal type_cast_1102_inst_req_1 : boolean;
  signal type_cast_1102_inst_ack_1 : boolean;
  signal if_stmt_1140_branch_req_0 : boolean;
  signal if_stmt_1140_branch_ack_1 : boolean;
  signal if_stmt_1140_branch_ack_0 : boolean;
  signal type_cast_1161_inst_req_0 : boolean;
  signal type_cast_1161_inst_ack_0 : boolean;
  signal type_cast_1161_inst_req_1 : boolean;
  signal type_cast_1161_inst_ack_1 : boolean;
  signal type_cast_1165_inst_req_0 : boolean;
  signal type_cast_1165_inst_ack_0 : boolean;
  signal type_cast_1165_inst_req_1 : boolean;
  signal type_cast_1165_inst_ack_1 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal type_cast_1174_inst_req_1 : boolean;
  signal type_cast_1174_inst_ack_1 : boolean;
  signal type_cast_1183_inst_req_0 : boolean;
  signal type_cast_1183_inst_ack_0 : boolean;
  signal type_cast_1183_inst_req_1 : boolean;
  signal type_cast_1183_inst_ack_1 : boolean;
  signal type_cast_1192_inst_req_0 : boolean;
  signal type_cast_1192_inst_ack_0 : boolean;
  signal type_cast_1192_inst_req_1 : boolean;
  signal type_cast_1192_inst_ack_1 : boolean;
  signal type_cast_1197_inst_req_0 : boolean;
  signal type_cast_1197_inst_ack_0 : boolean;
  signal type_cast_1197_inst_req_1 : boolean;
  signal type_cast_1197_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1357_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1357_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1357_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1357_inst_ack_1 : boolean;
  signal type_cast_1361_inst_req_0 : boolean;
  signal type_cast_1361_inst_ack_0 : boolean;
  signal type_cast_1361_inst_req_1 : boolean;
  signal type_cast_1361_inst_ack_1 : boolean;
  signal ptr_deref_1369_store_0_req_0 : boolean;
  signal ptr_deref_1369_store_0_ack_0 : boolean;
  signal ptr_deref_1369_store_0_req_1 : boolean;
  signal ptr_deref_1369_store_0_ack_1 : boolean;
  signal if_stmt_1383_branch_req_0 : boolean;
  signal if_stmt_1383_branch_ack_1 : boolean;
  signal if_stmt_1383_branch_ack_0 : boolean;
  signal if_stmt_1434_branch_req_0 : boolean;
  signal if_stmt_1434_branch_ack_1 : boolean;
  signal if_stmt_1434_branch_ack_0 : boolean;
  signal type_cast_1449_inst_req_0 : boolean;
  signal type_cast_754_inst_req_0 : boolean;
  signal type_cast_1449_inst_ack_0 : boolean;
  signal type_cast_1449_inst_req_1 : boolean;
  signal type_cast_1449_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1792_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1792_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1487_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1487_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1487_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1487_inst_ack_1 : boolean;
  signal phi_stmt_993_req_1 : boolean;
  signal type_cast_999_inst_ack_1 : boolean;
  signal type_cast_999_inst_req_1 : boolean;
  signal type_cast_1491_inst_req_0 : boolean;
  signal type_cast_1491_inst_ack_0 : boolean;
  signal type_cast_1491_inst_req_1 : boolean;
  signal type_cast_1491_inst_ack_1 : boolean;
  signal phi_stmt_945_req_1 : boolean;
  signal type_cast_1506_inst_req_0 : boolean;
  signal type_cast_1506_inst_ack_0 : boolean;
  signal type_cast_1506_inst_req_1 : boolean;
  signal type_cast_1506_inst_ack_1 : boolean;
  signal type_cast_1758_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1798_inst_ack_1 : boolean;
  signal if_stmt_1513_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1798_inst_req_1 : boolean;
  signal if_stmt_1513_branch_ack_1 : boolean;
  signal if_stmt_1513_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1780_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1798_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1789_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1789_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1798_inst_req_0 : boolean;
  signal phi_stmt_945_ack_0 : boolean;
  signal array_obj_ref_1552_index_offset_req_0 : boolean;
  signal array_obj_ref_1552_index_offset_ack_0 : boolean;
  signal array_obj_ref_1552_index_offset_req_1 : boolean;
  signal phi_stmt_751_req_1 : boolean;
  signal array_obj_ref_1552_index_offset_ack_1 : boolean;
  signal type_cast_999_inst_ack_0 : boolean;
  signal phi_stmt_993_req_0 : boolean;
  signal addr_of_1553_final_reg_req_0 : boolean;
  signal addr_of_1553_final_reg_ack_0 : boolean;
  signal addr_of_1553_final_reg_req_1 : boolean;
  signal addr_of_1553_final_reg_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1789_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1789_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1786_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1786_inst_req_1 : boolean;
  signal type_cast_1748_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1780_inst_req_1 : boolean;
  signal ptr_deref_1556_store_0_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1786_inst_ack_0 : boolean;
  signal ptr_deref_1556_store_0_ack_0 : boolean;
  signal ptr_deref_1556_store_0_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1786_inst_req_0 : boolean;
  signal ptr_deref_1556_store_0_ack_1 : boolean;
  signal type_cast_1768_inst_ack_1 : boolean;
  signal type_cast_1768_inst_req_1 : boolean;
  signal type_cast_999_inst_req_0 : boolean;
  signal call_stmt_1563_call_req_0 : boolean;
  signal call_stmt_1563_call_ack_0 : boolean;
  signal call_stmt_1563_call_req_1 : boolean;
  signal call_stmt_1563_call_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1575_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1575_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1575_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1575_inst_ack_1 : boolean;
  signal type_cast_1768_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1578_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1801_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1578_inst_ack_0 : boolean;
  signal type_cast_1768_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1578_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1801_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1578_inst_ack_1 : boolean;
  signal phi_stmt_945_req_0 : boolean;
  signal type_cast_948_inst_ack_1 : boolean;
  signal type_cast_948_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1582_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1783_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1783_inst_req_1 : boolean;
  signal type_cast_1606_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1801_inst_ack_0 : boolean;
  signal type_cast_1606_inst_ack_0 : boolean;
  signal type_cast_1606_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1801_inst_req_0 : boolean;
  signal type_cast_1606_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1783_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1783_inst_req_0 : boolean;
  signal type_cast_1616_inst_req_0 : boolean;
  signal type_cast_1616_inst_ack_0 : boolean;
  signal phi_stmt_986_req_0 : boolean;
  signal type_cast_1616_inst_req_1 : boolean;
  signal type_cast_1616_inst_ack_1 : boolean;
  signal type_cast_1625_inst_req_0 : boolean;
  signal type_cast_1625_inst_ack_0 : boolean;
  signal type_cast_1625_inst_req_1 : boolean;
  signal type_cast_1625_inst_ack_1 : boolean;
  signal type_cast_1654_inst_req_0 : boolean;
  signal type_cast_1654_inst_ack_0 : boolean;
  signal type_cast_1654_inst_req_1 : boolean;
  signal type_cast_1654_inst_ack_1 : boolean;
  signal type_cast_1658_inst_req_0 : boolean;
  signal type_cast_1658_inst_ack_0 : boolean;
  signal type_cast_1658_inst_req_1 : boolean;
  signal type_cast_1658_inst_ack_1 : boolean;
  signal call_stmt_1662_call_req_0 : boolean;
  signal call_stmt_1662_call_ack_0 : boolean;
  signal call_stmt_1662_call_req_1 : boolean;
  signal call_stmt_1662_call_ack_1 : boolean;
  signal call_stmt_1669_call_req_0 : boolean;
  signal call_stmt_1669_call_ack_0 : boolean;
  signal call_stmt_1669_call_req_1 : boolean;
  signal call_stmt_1669_call_ack_1 : boolean;
  signal if_stmt_1681_branch_req_0 : boolean;
  signal if_stmt_1681_branch_ack_1 : boolean;
  signal if_stmt_1681_branch_ack_0 : boolean;
  signal type_cast_1691_inst_req_0 : boolean;
  signal type_cast_1691_inst_ack_0 : boolean;
  signal type_cast_1691_inst_req_1 : boolean;
  signal type_cast_1691_inst_ack_1 : boolean;
  signal call_stmt_1695_call_req_0 : boolean;
  signal call_stmt_1695_call_ack_0 : boolean;
  signal call_stmt_1695_call_req_1 : boolean;
  signal call_stmt_1695_call_ack_1 : boolean;
  signal type_cast_1699_inst_req_0 : boolean;
  signal type_cast_1699_inst_ack_0 : boolean;
  signal type_cast_1699_inst_req_1 : boolean;
  signal type_cast_1699_inst_ack_1 : boolean;
  signal type_cast_1708_inst_req_0 : boolean;
  signal type_cast_1708_inst_ack_0 : boolean;
  signal type_cast_1708_inst_req_1 : boolean;
  signal type_cast_1708_inst_ack_1 : boolean;
  signal type_cast_1718_inst_req_0 : boolean;
  signal type_cast_1718_inst_ack_0 : boolean;
  signal type_cast_1718_inst_req_1 : boolean;
  signal type_cast_1718_inst_ack_1 : boolean;
  signal type_cast_1728_inst_req_0 : boolean;
  signal type_cast_1728_inst_ack_0 : boolean;
  signal type_cast_1728_inst_req_1 : boolean;
  signal type_cast_1728_inst_ack_1 : boolean;
  signal type_cast_1738_inst_req_0 : boolean;
  signal type_cast_1738_inst_ack_0 : boolean;
  signal type_cast_1738_inst_req_1 : boolean;
  signal type_cast_1738_inst_ack_1 : boolean;
  signal type_cast_1050_inst_req_0 : boolean;
  signal type_cast_1050_inst_ack_0 : boolean;
  signal type_cast_1050_inst_req_1 : boolean;
  signal type_cast_1050_inst_ack_1 : boolean;
  signal phi_stmt_1047_req_0 : boolean;
  signal phi_stmt_1047_ack_0 : boolean;
  signal phi_stmt_1220_req_0 : boolean;
  signal type_cast_1226_inst_req_0 : boolean;
  signal type_cast_1226_inst_ack_0 : boolean;
  signal type_cast_1226_inst_req_1 : boolean;
  signal type_cast_1226_inst_ack_1 : boolean;
  signal phi_stmt_1220_req_1 : boolean;
  signal phi_stmt_1220_ack_0 : boolean;
  signal type_cast_1417_inst_req_0 : boolean;
  signal type_cast_1417_inst_ack_0 : boolean;
  signal type_cast_1417_inst_req_1 : boolean;
  signal type_cast_1417_inst_ack_1 : boolean;
  signal phi_stmt_1414_req_0 : boolean;
  signal phi_stmt_1414_req_1 : boolean;
  signal phi_stmt_1414_ack_0 : boolean;
  signal phi_stmt_1459_req_0 : boolean;
  signal phi_stmt_1466_req_0 : boolean;
  signal type_cast_1465_inst_req_0 : boolean;
  signal type_cast_1465_inst_ack_0 : boolean;
  signal type_cast_1465_inst_req_1 : boolean;
  signal type_cast_1465_inst_ack_1 : boolean;
  signal phi_stmt_1459_req_1 : boolean;
  signal type_cast_1472_inst_req_0 : boolean;
  signal type_cast_1472_inst_ack_0 : boolean;
  signal type_cast_1472_inst_req_1 : boolean;
  signal type_cast_1472_inst_ack_1 : boolean;
  signal phi_stmt_1466_req_1 : boolean;
  signal phi_stmt_1459_ack_0 : boolean;
  signal phi_stmt_1466_ack_0 : boolean;
  signal type_cast_1523_inst_req_0 : boolean;
  signal type_cast_1523_inst_ack_0 : boolean;
  signal type_cast_1523_inst_req_1 : boolean;
  signal type_cast_1523_inst_ack_1 : boolean;
  signal phi_stmt_1520_req_0 : boolean;
  signal phi_stmt_1520_ack_0 : boolean;
  signal phi_stmt_1634_req_1 : boolean;
  signal type_cast_1637_inst_req_0 : boolean;
  signal type_cast_1637_inst_ack_0 : boolean;
  signal type_cast_1637_inst_req_1 : boolean;
  signal type_cast_1637_inst_ack_1 : boolean;
  signal phi_stmt_1634_req_0 : boolean;
  signal phi_stmt_1634_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_1115_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1115_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_1115_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_1115_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_1115: Block -- control-path 
    signal convolution3D_CP_1115_elements: BooleanArray(372 downto 0);
    -- 
  begin -- 
    convolution3D_CP_1115_elements(0) <= convolution3D_CP_1115_start;
    convolution3D_CP_1115_symbol <= convolution3D_CP_1115_elements(304);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	73 
    -- CP-element group 0:  members (65) 
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_441/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/branch_block_stmt_441__entry__
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672__entry__
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_update_start_
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Update/cr
      -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_586_inst_req_1); -- 
    cr_1530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_573_inst_req_1); -- 
    cr_1642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_623_inst_req_1); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_561_inst_req_1); -- 
    cr_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_548_inst_req_1); -- 
    cr_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_598_inst_req_1); -- 
    cr_1712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_665_inst_req_1); -- 
    cr_1698_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1698_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_649_inst_req_1); -- 
    cr_1670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_636_inst_req_1); -- 
    cr_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_611_inst_req_1); -- 
    cr_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_511_inst_req_1); -- 
    cr_1684_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1684_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_645_inst_req_1); -- 
    cr_1446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_536_inst_req_1); -- 
    cr_1418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_523_inst_req_1); -- 
    rr_1231_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1231_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => RPIPE_maxpool_input_pipe_444_inst_req_0); -- 
    cr_1250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_448_inst_req_1); -- 
    cr_1278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_461_inst_req_1); -- 
    cr_1306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_473_inst_req_1); -- 
    cr_1334_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1334_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_486_inst_req_1); -- 
    cr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(0), ack => type_cast_498_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_update_start_
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Update/cr
      -- 
    ra_1232_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_444_inst_ack_0, ack => convolution3D_CP_1115_elements(1)); -- 
    cr_1236_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1236_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(1), ack => RPIPE_maxpool_input_pipe_444_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_444_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Sample/rr
      -- 
    ca_1237_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_444_inst_ack_1, ack => convolution3D_CP_1115_elements(2)); -- 
    rr_1245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(2), ack => type_cast_448_inst_req_0); -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(2), ack => RPIPE_maxpool_input_pipe_457_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Sample/ra
      -- 
    ra_1246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_448_inst_ack_0, ack => convolution3D_CP_1115_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_448_Update/ca
      -- 
    ca_1251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_448_inst_ack_1, ack => convolution3D_CP_1115_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_update_start_
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Update/cr
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_457_inst_ack_0, ack => convolution3D_CP_1115_elements(5)); -- 
    cr_1264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(5), ack => RPIPE_maxpool_input_pipe_457_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_457_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Sample/rr
      -- 
    ca_1265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_457_inst_ack_1, ack => convolution3D_CP_1115_elements(6)); -- 
    rr_1273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(6), ack => type_cast_461_inst_req_0); -- 
    rr_1287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(6), ack => RPIPE_maxpool_input_pipe_469_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Sample/ra
      -- 
    ra_1274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_0, ack => convolution3D_CP_1115_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_461_Update/ca
      -- 
    ca_1279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_461_inst_ack_1, ack => convolution3D_CP_1115_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_update_start_
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Update/cr
      -- 
    ra_1288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_0, ack => convolution3D_CP_1115_elements(9)); -- 
    cr_1292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(9), ack => RPIPE_maxpool_input_pipe_469_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_469_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Sample/rr
      -- 
    ca_1293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_469_inst_ack_1, ack => convolution3D_CP_1115_elements(10)); -- 
    rr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1301_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(10), ack => type_cast_473_inst_req_0); -- 
    rr_1315_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1315_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(10), ack => RPIPE_maxpool_input_pipe_482_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Sample/ra
      -- 
    ra_1302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_0, ack => convolution3D_CP_1115_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_473_Update/ca
      -- 
    ca_1307_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_473_inst_ack_1, ack => convolution3D_CP_1115_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_update_start_
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Update/cr
      -- 
    ra_1316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_482_inst_ack_0, ack => convolution3D_CP_1115_elements(13)); -- 
    cr_1320_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1320_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(13), ack => RPIPE_maxpool_input_pipe_482_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_482_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Sample/rr
      -- 
    ca_1321_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_482_inst_ack_1, ack => convolution3D_CP_1115_elements(14)); -- 
    rr_1329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(14), ack => type_cast_486_inst_req_0); -- 
    rr_1343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(14), ack => RPIPE_maxpool_input_pipe_494_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Sample/ra
      -- 
    ra_1330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => convolution3D_CP_1115_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_486_Update/ca
      -- 
    ca_1335_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => convolution3D_CP_1115_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_update_start_
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Update/cr
      -- 
    ra_1344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_494_inst_ack_0, ack => convolution3D_CP_1115_elements(17)); -- 
    cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(17), ack => RPIPE_maxpool_input_pipe_494_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_494_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_sample_start_
      -- 
    ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_494_inst_ack_1, ack => convolution3D_CP_1115_elements(18)); -- 
    rr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(18), ack => type_cast_498_inst_req_0); -- 
    rr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(18), ack => RPIPE_maxpool_input_pipe_507_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Sample/ra
      -- 
    ra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_0, ack => convolution3D_CP_1115_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_498_Update/ca
      -- 
    ca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_498_inst_ack_1, ack => convolution3D_CP_1115_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Update/$entry
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_update_start_
      -- 
    ra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_507_inst_ack_0, ack => convolution3D_CP_1115_elements(21)); -- 
    cr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(21), ack => RPIPE_maxpool_input_pipe_507_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22: 	25 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_507_update_completed_
      -- 
    ca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_507_inst_ack_1, ack => convolution3D_CP_1115_elements(22)); -- 
    rr_1385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(22), ack => type_cast_511_inst_req_0); -- 
    rr_1399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(22), ack => RPIPE_maxpool_input_pipe_519_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Sample/ra
      -- 
    ra_1386_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_0, ack => convolution3D_CP_1115_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_511_Update/ca
      -- 
    ca_1391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_511_inst_ack_1, ack => convolution3D_CP_1115_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_update_start_
      -- CP-element group 25: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_sample_completed_
      -- 
    ra_1400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_519_inst_ack_0, ack => convolution3D_CP_1115_elements(25)); -- 
    cr_1404_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1404_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(25), ack => RPIPE_maxpool_input_pipe_519_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_519_update_completed_
      -- 
    ca_1405_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_519_inst_ack_1, ack => convolution3D_CP_1115_elements(26)); -- 
    rr_1413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(26), ack => type_cast_523_inst_req_0); -- 
    rr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(26), ack => RPIPE_maxpool_input_pipe_532_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Sample/ra
      -- 
    ra_1414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_0, ack => convolution3D_CP_1115_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	74 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_523_Update/$exit
      -- 
    ca_1419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_523_inst_ack_1, ack => convolution3D_CP_1115_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Sample/ra
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_update_start_
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_sample_completed_
      -- 
    ra_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_532_inst_ack_0, ack => convolution3D_CP_1115_elements(29)); -- 
    cr_1432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(29), ack => RPIPE_maxpool_input_pipe_532_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_532_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Sample/rr
      -- 
    ca_1433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_532_inst_ack_1, ack => convolution3D_CP_1115_elements(30)); -- 
    rr_1441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(30), ack => type_cast_536_inst_req_0); -- 
    rr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(30), ack => RPIPE_maxpool_input_pipe_544_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Sample/ra
      -- 
    ra_1442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_0, ack => convolution3D_CP_1115_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	74 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_536_Update/ca
      -- 
    ca_1447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_536_inst_ack_1, ack => convolution3D_CP_1115_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_update_start_
      -- CP-element group 33: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Sample/ra
      -- 
    ra_1456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_544_inst_ack_0, ack => convolution3D_CP_1115_elements(33)); -- 
    cr_1460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(33), ack => RPIPE_maxpool_input_pipe_544_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	37 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_544_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Sample/$entry
      -- 
    ca_1461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_544_inst_ack_1, ack => convolution3D_CP_1115_elements(34)); -- 
    rr_1469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(34), ack => type_cast_548_inst_req_0); -- 
    rr_1483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(34), ack => RPIPE_maxpool_input_pipe_557_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_sample_completed_
      -- 
    ra_1470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_0, ack => convolution3D_CP_1115_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	74 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_548_update_completed_
      -- 
    ca_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_1, ack => convolution3D_CP_1115_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_update_start_
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Sample/$exit
      -- 
    ra_1484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_0, ack => convolution3D_CP_1115_elements(37)); -- 
    cr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(37), ack => RPIPE_maxpool_input_pipe_557_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_557_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_sample_start_
      -- 
    ca_1489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_557_inst_ack_1, ack => convolution3D_CP_1115_elements(38)); -- 
    rr_1497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(38), ack => type_cast_561_inst_req_0); -- 
    rr_1511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(38), ack => RPIPE_maxpool_input_pipe_569_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Sample/ra
      -- 
    ra_1498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => convolution3D_CP_1115_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	74 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_561_Update/ca
      -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => convolution3D_CP_1115_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Update/cr
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_update_start_
      -- CP-element group 41: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_sample_completed_
      -- 
    ra_1512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_569_inst_ack_0, ack => convolution3D_CP_1115_elements(41)); -- 
    cr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(41), ack => RPIPE_maxpool_input_pipe_569_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_569_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Sample/$entry
      -- 
    ca_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_569_inst_ack_1, ack => convolution3D_CP_1115_elements(42)); -- 
    rr_1525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(42), ack => type_cast_573_inst_req_0); -- 
    rr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(42), ack => RPIPE_maxpool_input_pipe_582_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Sample/$exit
      -- 
    ra_1526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => convolution3D_CP_1115_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	74 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_573_Update/ca
      -- 
    ca_1531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_1, ack => convolution3D_CP_1115_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_update_start_
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Update/cr
      -- 
    ra_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_0, ack => convolution3D_CP_1115_elements(45)); -- 
    cr_1544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(45), ack => RPIPE_maxpool_input_pipe_582_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_582_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Sample/rr
      -- 
    ca_1545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_582_inst_ack_1, ack => convolution3D_CP_1115_elements(46)); -- 
    rr_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(46), ack => type_cast_586_inst_req_0); -- 
    rr_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(46), ack => RPIPE_maxpool_input_pipe_594_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Sample/$exit
      -- 
    ra_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_0, ack => convolution3D_CP_1115_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	74 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_586_Update/ca
      -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_586_inst_ack_1, ack => convolution3D_CP_1115_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_update_start_
      -- 
    ra_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_594_inst_ack_0, ack => convolution3D_CP_1115_elements(49)); -- 
    cr_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(49), ack => RPIPE_maxpool_input_pipe_594_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_594_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Sample/$entry
      -- 
    ca_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_594_inst_ack_1, ack => convolution3D_CP_1115_elements(50)); -- 
    rr_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(50), ack => type_cast_598_inst_req_0); -- 
    rr_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(50), ack => RPIPE_maxpool_input_pipe_607_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Sample/ra
      -- 
    ra_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_0, ack => convolution3D_CP_1115_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	74 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_598_update_completed_
      -- 
    ca_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_598_inst_ack_1, ack => convolution3D_CP_1115_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_update_start_
      -- 
    ra_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_0, ack => convolution3D_CP_1115_elements(53)); -- 
    cr_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(53), ack => RPIPE_maxpool_input_pipe_607_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_607_update_completed_
      -- 
    ca_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_607_inst_ack_1, ack => convolution3D_CP_1115_elements(54)); -- 
    rr_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(54), ack => type_cast_611_inst_req_0); -- 
    rr_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(54), ack => RPIPE_maxpool_input_pipe_619_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Sample/$exit
      -- 
    ra_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_0, ack => convolution3D_CP_1115_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	74 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_611_update_completed_
      -- 
    ca_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_611_inst_ack_1, ack => convolution3D_CP_1115_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Update/cr
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_update_start_
      -- 
    ra_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_619_inst_ack_0, ack => convolution3D_CP_1115_elements(57)); -- 
    cr_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(57), ack => RPIPE_maxpool_input_pipe_619_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	61 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_619_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Sample/rr
      -- 
    ca_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_619_inst_ack_1, ack => convolution3D_CP_1115_elements(58)); -- 
    rr_1637_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1637_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(58), ack => type_cast_623_inst_req_0); -- 
    rr_1651_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1651_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(58), ack => RPIPE_maxpool_input_pipe_632_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Sample/ra
      -- CP-element group 59: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Sample/$exit
      -- 
    ra_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_0, ack => convolution3D_CP_1115_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	74 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_623_Update/$exit
      -- 
    ca_1643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_623_inst_ack_1, ack => convolution3D_CP_1115_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_update_start_
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Update/cr
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Sample/$exit
      -- 
    ra_1652_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_0, ack => convolution3D_CP_1115_elements(61)); -- 
    cr_1656_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1656_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(61), ack => RPIPE_maxpool_input_pipe_632_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/RPIPE_maxpool_input_pipe_632_Update/$exit
      -- 
    ca_1657_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_632_inst_ack_1, ack => convolution3D_CP_1115_elements(62)); -- 
    rr_1665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(62), ack => type_cast_636_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_sample_completed_
      -- 
    ra_1666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => convolution3D_CP_1115_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	74 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_636_update_completed_
      -- 
    ca_1671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_1, ack => convolution3D_CP_1115_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	16 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Sample/$entry
      -- 
    rr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(65), ack => type_cast_645_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(12) & convolution3D_CP_1115_elements(16);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_sample_completed_
      -- 
    ra_1680_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_0, ack => convolution3D_CP_1115_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_645_Update/$exit
      -- 
    ca_1685_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_645_inst_ack_1, ack => convolution3D_CP_1115_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_sample_start_
      -- 
    rr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(68), ack => type_cast_649_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(20) & convolution3D_CP_1115_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Sample/ra
      -- CP-element group 69: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_sample_completed_
      -- 
    ra_1694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => convolution3D_CP_1115_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_649_Update/ca
      -- 
    ca_1699_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => convolution3D_CP_1115_elements(70)); -- 
    -- CP-element group 71:  join  transition  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Sample/rr
      -- 
    rr_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(71), ack => type_cast_665_inst_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(4) & convolution3D_CP_1115_elements(8) & convolution3D_CP_1115_elements(67) & convolution3D_CP_1115_elements(70);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Sample/$exit
      -- 
    ra_1708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_0, ack => convolution3D_CP_1115_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	0 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/type_cast_665_Update/$exit
      -- 
    ca_1713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_1, ack => convolution3D_CP_1115_elements(73)); -- 
    -- CP-element group 74:  branch  join  transition  place  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: 	32 
    -- CP-element group 74: 	36 
    -- CP-element group 74: 	40 
    -- CP-element group 74: 	44 
    -- CP-element group 74: 	48 
    -- CP-element group 74: 	52 
    -- CP-element group 74: 	56 
    -- CP-element group 74: 	60 
    -- CP-element group 74: 	64 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (10) 
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_else_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_eval_test/$exit
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_if_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_eval_test/branch_req
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_eval_test/$entry
      -- CP-element group 74: 	 branch_block_stmt_441/R_cmp383_674_place
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673_dead_link/$entry
      -- CP-element group 74: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672__exit__
      -- CP-element group 74: 	 branch_block_stmt_441/if_stmt_673__entry__
      -- CP-element group 74: 	 branch_block_stmt_441/assign_stmt_445_to_assign_stmt_672/$exit
      -- 
    branch_req_1721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(74), ack => if_stmt_673_branch_req_0); -- 
    convolution3D_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(28) & convolution3D_CP_1115_elements(32) & convolution3D_CP_1115_elements(36) & convolution3D_CP_1115_elements(40) & convolution3D_CP_1115_elements(44) & convolution3D_CP_1115_elements(48) & convolution3D_CP_1115_elements(52) & convolution3D_CP_1115_elements(56) & convolution3D_CP_1115_elements(60) & convolution3D_CP_1115_elements(64) & convolution3D_CP_1115_elements(73);
      gj_convolution3D_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: 	78 
    -- CP-element group 75: 	79 
    -- CP-element group 75: 	80 
    -- CP-element group 75: 	81 
    -- CP-element group 75: 	82 
    -- CP-element group 75: 	85 
    -- CP-element group 75:  members (33) 
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_update_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_update_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_update_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Sample/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/if_stmt_673_if_link/if_choice_transition
      -- CP-element group 75: 	 branch_block_stmt_441/if_stmt_673_if_link/$exit
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_update_start_
      -- CP-element group 75: 	 branch_block_stmt_441/entry_bbx_xnph385
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_441/merge_stmt_679__exit__
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748__entry__
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Update/cr
      -- CP-element group 75: 	 branch_block_stmt_441/merge_stmt_679_PhiAck/dummy
      -- CP-element group 75: 	 branch_block_stmt_441/merge_stmt_679_PhiAck/$exit
      -- CP-element group 75: 	 branch_block_stmt_441/merge_stmt_679_PhiAck/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/entry_bbx_xnph385_PhiReq/$exit
      -- CP-element group 75: 	 branch_block_stmt_441/entry_bbx_xnph385_PhiReq/$entry
      -- CP-element group 75: 	 branch_block_stmt_441/merge_stmt_679_PhiReqMerge
      -- 
    if_choice_transition_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_673_branch_ack_1, ack => convolution3D_CP_1115_elements(75)); -- 
    rr_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_718_inst_req_0); -- 
    cr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_693_inst_req_1); -- 
    rr_1743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_693_inst_req_0); -- 
    rr_1757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_709_inst_req_0); -- 
    cr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_709_inst_req_1); -- 
    cr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_718_inst_req_1); -- 
    cr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(75), ack => type_cast_728_inst_req_1); -- 
    -- CP-element group 76:  transition  place  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	311 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_441/if_stmt_673_else_link/else_choice_transition
      -- CP-element group 76: 	 branch_block_stmt_441/if_stmt_673_else_link/$exit
      -- CP-element group 76: 	 branch_block_stmt_441/entry_forx_xend
      -- CP-element group 76: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/$entry
      -- CP-element group 76: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/$entry
      -- CP-element group 76: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_1730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_673_branch_ack_0, ack => convolution3D_CP_1115_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_sample_completed_
      -- 
    ra_1744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_0, ack => convolution3D_CP_1115_elements(77)); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	75 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	86 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_693_Update/ca
      -- 
    ca_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_693_inst_ack_1, ack => convolution3D_CP_1115_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	75 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Sample/ra
      -- 
    ra_1758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_0, ack => convolution3D_CP_1115_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	75 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	83 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_709_Update/ca
      -- 
    ca_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_709_inst_ack_1, ack => convolution3D_CP_1115_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	75 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Sample/ra
      -- 
    ra_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_0, ack => convolution3D_CP_1115_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	75 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_718_Update/ca
      -- 
    ca_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_718_inst_ack_1, ack => convolution3D_CP_1115_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	80 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Sample/rr
      -- 
    rr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(83), ack => type_cast_728_inst_req_0); -- 
    convolution3D_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(80) & convolution3D_CP_1115_elements(82);
      gj_convolution3D_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Sample/ra
      -- 
    ra_1786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_0, ack => convolution3D_CP_1115_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	75 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/type_cast_728_Update/ca
      -- 
    ca_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_728_inst_ack_1, ack => convolution3D_CP_1115_elements(85)); -- 
    -- CP-element group 86:  join  transition  place  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	78 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	305 
    -- CP-element group 86:  members (6) 
      -- CP-element group 86: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748/$exit
      -- CP-element group 86: 	 branch_block_stmt_441/assign_stmt_684_to_assign_stmt_748__exit__
      -- CP-element group 86: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody
      -- CP-element group 86: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/$entry
      -- CP-element group 86: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/$entry
      -- CP-element group 86: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(78) & convolution3D_CP_1115_elements(85);
      gj_convolution3D_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	310 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	126 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_sample_complete
      -- CP-element group 87: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Sample/ack
      -- 
    ack_1820_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_763_index_offset_ack_0, ack => convolution3D_CP_1115_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	310 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (11) 
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_root_address_calculated
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_offset_calculated
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Update/ack
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_base_plus_offset/$entry
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_base_plus_offset/$exit
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_base_plus_offset/sum_rename_req
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_base_plus_offset/sum_rename_ack
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_request/$entry
      -- CP-element group 88: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_request/req
      -- 
    ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_763_index_offset_ack_1, ack => convolution3D_CP_1115_elements(88)); -- 
    req_1834_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1834_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(88), ack => addr_of_764_final_reg_req_0); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_request/$exit
      -- CP-element group 89: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_request/ack
      -- 
    ack_1835_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_764_final_reg_ack_0, ack => convolution3D_CP_1115_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	310 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	123 
    -- CP-element group 90:  members (19) 
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_complete/$exit
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_complete/ack
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_word_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_root_address_calculated
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_address_resized
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_addr_resize/$entry
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_addr_resize/$exit
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_addr_resize/base_resize_req
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_addr_resize/base_resize_ack
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_plus_offset/$entry
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_plus_offset/$exit
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_plus_offset/sum_rename_req
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_base_plus_offset/sum_rename_ack
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_word_addrgen/$entry
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_word_addrgen/$exit
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_word_addrgen/root_register_req
      -- CP-element group 90: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_word_addrgen/root_register_ack
      -- 
    ack_1840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_764_final_reg_ack_1, ack => convolution3D_CP_1115_elements(90)); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	310 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_update_start_
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Update/cr
      -- 
    ra_1849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_767_inst_ack_0, ack => convolution3D_CP_1115_elements(91)); -- 
    cr_1853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(91), ack => RPIPE_maxpool_input_pipe_767_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92: 	95 
    -- CP-element group 92:  members (9) 
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Update/$exit
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Update/ca
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Sample/rr
      -- 
    ca_1854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_767_inst_ack_1, ack => convolution3D_CP_1115_elements(92)); -- 
    rr_1862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(92), ack => type_cast_771_inst_req_0); -- 
    rr_1876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(92), ack => RPIPE_maxpool_input_pipe_780_inst_req_0); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Sample/ra
      -- 
    ra_1863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_771_inst_ack_0, ack => convolution3D_CP_1115_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	310 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	123 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Update/ca
      -- 
    ca_1868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_771_inst_ack_1, ack => convolution3D_CP_1115_elements(94)); -- 
    -- CP-element group 95:  transition  input  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	92 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_update_start_
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Update/$entry
      -- CP-element group 95: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Update/cr
      -- 
    ra_1877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_780_inst_ack_0, ack => convolution3D_CP_1115_elements(95)); -- 
    cr_1881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(95), ack => RPIPE_maxpool_input_pipe_780_inst_req_1); -- 
    -- CP-element group 96:  fork  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	95 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96: 	99 
    -- CP-element group 96:  members (9) 
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_update_completed_
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_780_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Sample/rr
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Sample/rr
      -- 
    ca_1882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_780_inst_ack_1, ack => convolution3D_CP_1115_elements(96)); -- 
    rr_1890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(96), ack => type_cast_784_inst_req_0); -- 
    rr_1904_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1904_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(96), ack => RPIPE_maxpool_input_pipe_798_inst_req_0); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Sample/ra
      -- 
    ra_1891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_0, ack => convolution3D_CP_1115_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	310 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	123 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Update/ca
      -- 
    ca_1896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_784_inst_ack_1, ack => convolution3D_CP_1115_elements(98)); -- 
    -- CP-element group 99:  transition  input  output  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	96 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (6) 
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_update_start_
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Update/$entry
      -- CP-element group 99: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Update/cr
      -- 
    ra_1905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_798_inst_ack_0, ack => convolution3D_CP_1115_elements(99)); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1909_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(99), ack => RPIPE_maxpool_input_pipe_798_inst_req_1); -- 
    -- CP-element group 100:  fork  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_798_Update/ca
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Sample/rr
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_sample_start_
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Sample/$entry
      -- CP-element group 100: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Sample/rr
      -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_798_inst_ack_1, ack => convolution3D_CP_1115_elements(100)); -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(100), ack => type_cast_802_inst_req_0); -- 
    rr_1932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(100), ack => RPIPE_maxpool_input_pipe_816_inst_req_0); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Sample/ra
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_802_inst_ack_0, ack => convolution3D_CP_1115_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	310 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	123 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Update/ca
      -- 
    ca_1924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_802_inst_ack_1, ack => convolution3D_CP_1115_elements(102)); -- 
    -- CP-element group 103:  transition  input  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	100 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (6) 
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_update_start_
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Sample/ra
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Update/cr
      -- 
    ra_1933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_816_inst_ack_0, ack => convolution3D_CP_1115_elements(103)); -- 
    cr_1937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(103), ack => RPIPE_maxpool_input_pipe_816_inst_req_1); -- 
    -- CP-element group 104:  fork  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	107 
    -- CP-element group 104:  members (9) 
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_816_Update/ca
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Sample/rr
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Sample/rr
      -- 
    ca_1938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_816_inst_ack_1, ack => convolution3D_CP_1115_elements(104)); -- 
    rr_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(104), ack => type_cast_820_inst_req_0); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(104), ack => RPIPE_maxpool_input_pipe_834_inst_req_0); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Sample/ra
      -- 
    ra_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_820_inst_ack_0, ack => convolution3D_CP_1115_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	310 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	123 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Update/ca
      -- 
    ca_1952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_820_inst_ack_1, ack => convolution3D_CP_1115_elements(106)); -- 
    -- CP-element group 107:  transition  input  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	104 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (6) 
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_sample_completed_
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_update_start_
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Update/cr
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_834_inst_ack_0, ack => convolution3D_CP_1115_elements(107)); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(107), ack => RPIPE_maxpool_input_pipe_834_inst_req_1); -- 
    -- CP-element group 108:  fork  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108: 	111 
    -- CP-element group 108:  members (9) 
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_834_Update/ca
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Sample/rr
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Sample/rr
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_834_inst_ack_1, ack => convolution3D_CP_1115_elements(108)); -- 
    rr_1974_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1974_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(108), ack => type_cast_838_inst_req_0); -- 
    rr_1988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(108), ack => RPIPE_maxpool_input_pipe_852_inst_req_0); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Sample/ra
      -- 
    ra_1975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_0, ack => convolution3D_CP_1115_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	310 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	123 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Update/ca
      -- 
    ca_1980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_838_inst_ack_1, ack => convolution3D_CP_1115_elements(110)); -- 
    -- CP-element group 111:  transition  input  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	108 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (6) 
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_sample_completed_
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_update_start_
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Sample/$exit
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Sample/ra
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Update/cr
      -- 
    ra_1989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_852_inst_ack_0, ack => convolution3D_CP_1115_elements(111)); -- 
    cr_1993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(111), ack => RPIPE_maxpool_input_pipe_852_inst_req_1); -- 
    -- CP-element group 112:  fork  transition  input  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112: 	115 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_update_completed_
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Update/$exit
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_852_Update/ca
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Sample/rr
      -- 
    ca_1994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_852_inst_ack_1, ack => convolution3D_CP_1115_elements(112)); -- 
    rr_2002_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2002_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(112), ack => type_cast_856_inst_req_0); -- 
    rr_2016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(112), ack => RPIPE_maxpool_input_pipe_870_inst_req_0); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Sample/ra
      -- 
    ra_2003_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_0, ack => convolution3D_CP_1115_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	310 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	123 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Update/ca
      -- 
    ca_2008_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_856_inst_ack_1, ack => convolution3D_CP_1115_elements(114)); -- 
    -- CP-element group 115:  transition  input  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	112 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_update_start_
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Update/cr
      -- 
    ra_2017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_870_inst_ack_0, ack => convolution3D_CP_1115_elements(115)); -- 
    cr_2021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(115), ack => RPIPE_maxpool_input_pipe_870_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (9) 
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_870_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Sample/rr
      -- 
    ca_2022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_870_inst_ack_1, ack => convolution3D_CP_1115_elements(116)); -- 
    rr_2030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(116), ack => type_cast_874_inst_req_0); -- 
    rr_2044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(116), ack => RPIPE_maxpool_input_pipe_888_inst_req_0); -- 
    -- CP-element group 117:  transition  input  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	116 
    -- CP-element group 117: successors 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Sample/ra
      -- 
    ra_2031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_0, ack => convolution3D_CP_1115_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	310 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	123 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Update/ca
      -- 
    ca_2036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_874_inst_ack_1, ack => convolution3D_CP_1115_elements(118)); -- 
    -- CP-element group 119:  transition  input  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (6) 
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_update_start_
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Sample/ra
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Update/cr
      -- 
    ra_2045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_888_inst_ack_0, ack => convolution3D_CP_1115_elements(119)); -- 
    cr_2049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(119), ack => RPIPE_maxpool_input_pipe_888_inst_req_1); -- 
    -- CP-element group 120:  transition  input  output  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (6) 
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_888_Update/ca
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Sample/rr
      -- 
    ca_2050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_888_inst_ack_1, ack => convolution3D_CP_1115_elements(120)); -- 
    rr_2058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(120), ack => type_cast_892_inst_req_0); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Sample/ra
      -- 
    ra_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_892_inst_ack_0, ack => convolution3D_CP_1115_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	310 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Update/ca
      -- 
    ca_2064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_892_inst_ack_1, ack => convolution3D_CP_1115_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	90 
    -- CP-element group 123: 	94 
    -- CP-element group 123: 	98 
    -- CP-element group 123: 	102 
    -- CP-element group 123: 	106 
    -- CP-element group 123: 	110 
    -- CP-element group 123: 	114 
    -- CP-element group 123: 	118 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	124 
    -- CP-element group 123:  members (9) 
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/ptr_deref_900_Split/$entry
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/ptr_deref_900_Split/$exit
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/ptr_deref_900_Split/split_req
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/ptr_deref_900_Split/split_ack
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/$entry
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/word_0/$entry
      -- CP-element group 123: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/word_0/rr
      -- 
    rr_2102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(123), ack => ptr_deref_900_store_0_req_0); -- 
    convolution3D_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(90) & convolution3D_CP_1115_elements(94) & convolution3D_CP_1115_elements(98) & convolution3D_CP_1115_elements(102) & convolution3D_CP_1115_elements(106) & convolution3D_CP_1115_elements(110) & convolution3D_CP_1115_elements(114) & convolution3D_CP_1115_elements(118) & convolution3D_CP_1115_elements(122);
      gj_convolution3D_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	123 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (5) 
      -- CP-element group 124: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/$exit
      -- CP-element group 124: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/word_0/$exit
      -- CP-element group 124: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Sample/word_access_start/word_0/ra
      -- 
    ra_2103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_900_store_0_ack_0, ack => convolution3D_CP_1115_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	310 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	126 
    -- CP-element group 125:  members (5) 
      -- CP-element group 125: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/$exit
      -- CP-element group 125: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/word_0/$exit
      -- CP-element group 125: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/word_0/ca
      -- 
    ca_2114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_900_store_0_ack_1, ack => convolution3D_CP_1115_elements(125)); -- 
    -- CP-element group 126:  branch  join  transition  place  output  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	87 
    -- CP-element group 126: 	125 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	127 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (10) 
      -- CP-element group 126: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913__exit__
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914__entry__
      -- CP-element group 126: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/$exit
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_dead_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_eval_test/$entry
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_eval_test/$exit
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_eval_test/branch_req
      -- CP-element group 126: 	 branch_block_stmt_441/R_exitcond32_915_place
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_if_link/$entry
      -- CP-element group 126: 	 branch_block_stmt_441/if_stmt_914_else_link/$entry
      -- 
    branch_req_2122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(126), ack => if_stmt_914_branch_req_0); -- 
    convolution3D_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(87) & convolution3D_CP_1115_elements(125);
      gj_convolution3D_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	126 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	312 
    -- CP-element group 127: 	313 
    -- CP-element group 127:  members (24) 
      -- CP-element group 127: 	 branch_block_stmt_441/merge_stmt_920__exit__
      -- CP-element group 127: 	 branch_block_stmt_441/assign_stmt_927_to_assign_stmt_942__entry__
      -- CP-element group 127: 	 branch_block_stmt_441/assign_stmt_927_to_assign_stmt_942__exit__
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/rr
      -- CP-element group 127: 	 branch_block_stmt_441/if_stmt_914_if_link/$exit
      -- CP-element group 127: 	 branch_block_stmt_441/if_stmt_914_if_link/if_choice_transition
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xbody_forx_xcondx_xforx_xend_crit_edge
      -- CP-element group 127: 	 branch_block_stmt_441/assign_stmt_927_to_assign_stmt_942/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/assign_stmt_927_to_assign_stmt_942/$exit
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/merge_stmt_920_PhiAck/dummy
      -- CP-element group 127: 	 branch_block_stmt_441/merge_stmt_920_PhiReqMerge
      -- CP-element group 127: 	 branch_block_stmt_441/merge_stmt_920_PhiAck/$exit
      -- CP-element group 127: 	 branch_block_stmt_441/merge_stmt_920_PhiAck/$entry
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/cr
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$exit
      -- CP-element group 127: 	 branch_block_stmt_441/forx_xbody_forx_xcondx_xforx_xend_crit_edge_PhiReq/$entry
      -- 
    if_choice_transition_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_914_branch_ack_1, ack => convolution3D_CP_1115_elements(127)); -- 
    rr_3586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(127), ack => type_cast_948_inst_req_0); -- 
    cr_3591_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3591_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(127), ack => type_cast_948_inst_req_1); -- 
    -- CP-element group 128:  fork  transition  place  input  output  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	306 
    -- CP-element group 128: 	307 
    -- CP-element group 128:  members (12) 
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/cr
      -- CP-element group 128: 	 branch_block_stmt_441/if_stmt_914_else_link/$exit
      -- CP-element group 128: 	 branch_block_stmt_441/if_stmt_914_else_link/else_choice_transition
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/rr
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/$entry
      -- CP-element group 128: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_2131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_914_branch_ack_0, ack => convolution3D_CP_1115_elements(128)); -- 
    cr_3537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(128), ack => type_cast_754_inst_req_1); -- 
    rr_3532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(128), ack => type_cast_754_inst_req_0); -- 
    -- CP-element group 129:  transition  place  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	316 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	335 
    -- CP-element group 129:  members (5) 
      -- CP-element group 129: 	 branch_block_stmt_441/if_stmt_965_if_link/$exit
      -- CP-element group 129: 	 branch_block_stmt_441/if_stmt_965_if_link/if_choice_transition
      -- CP-element group 129: 	 branch_block_stmt_441/forx_xend_ifx_xend
      -- CP-element group 129: 	 branch_block_stmt_441/forx_xend_ifx_xend_PhiReq/$entry
      -- CP-element group 129: 	 branch_block_stmt_441/forx_xend_ifx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_1, ack => convolution3D_CP_1115_elements(129)); -- 
    -- CP-element group 130:  merge  fork  transition  place  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	316 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	317 
    -- CP-element group 130: 	318 
    -- CP-element group 130:  members (20) 
      -- CP-element group 130: 	 branch_block_stmt_441/merge_stmt_971__exit__
      -- CP-element group 130: 	 branch_block_stmt_441/assign_stmt_977_to_assign_stmt_983__entry__
      -- CP-element group 130: 	 branch_block_stmt_441/assign_stmt_977_to_assign_stmt_983__exit__
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi
      -- CP-element group 130: 	 branch_block_stmt_441/forx_xend_bbx_xnphx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/forx_xend_bbx_xnphx_xi_PhiReq/$exit
      -- CP-element group 130: 	 branch_block_stmt_441/merge_stmt_971_PhiAck/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/if_stmt_965_else_link/$exit
      -- CP-element group 130: 	 branch_block_stmt_441/if_stmt_965_else_link/else_choice_transition
      -- CP-element group 130: 	 branch_block_stmt_441/forx_xend_bbx_xnphx_xi
      -- CP-element group 130: 	 branch_block_stmt_441/assign_stmt_977_to_assign_stmt_983/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/assign_stmt_977_to_assign_stmt_983/$exit
      -- CP-element group 130: 	 branch_block_stmt_441/merge_stmt_971_PhiAck/$exit
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/merge_stmt_971_PhiReqMerge
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/merge_stmt_971_PhiAck/dummy
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/$entry
      -- CP-element group 130: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/$entry
      -- 
    else_choice_transition_2156_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_965_branch_ack_0, ack => convolution3D_CP_1115_elements(130)); -- 
    -- CP-element group 131:  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	330 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (6) 
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_sample_completed_
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_update_start_
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Sample/$exit
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Sample/ra
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Update/$entry
      -- CP-element group 131: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Update/cr
      -- 
    ra_2173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1014_inst_ack_0, ack => convolution3D_CP_1115_elements(131)); -- 
    cr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(131), ack => RPIPE_maxpool_input_pipe_1014_inst_req_1); -- 
    -- CP-element group 132:  transition  input  output  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	133 
    -- CP-element group 132:  members (6) 
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_update_completed_
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Update/ca
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Sample/rr
      -- 
    ca_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1014_inst_ack_1, ack => convolution3D_CP_1115_elements(132)); -- 
    rr_2186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(132), ack => type_cast_1018_inst_req_0); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	132 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Sample/ra
      -- 
    ra_2187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1018_inst_ack_0, ack => convolution3D_CP_1115_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	330 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	137 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Update/ca
      -- 
    ca_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1018_inst_ack_1, ack => convolution3D_CP_1115_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	330 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_sample_completed_
      -- CP-element group 135: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Sample/$exit
      -- CP-element group 135: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Sample/ra
      -- 
    ra_2201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_0, ack => convolution3D_CP_1115_elements(135)); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	330 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_update_completed_
      -- CP-element group 136: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Update/$exit
      -- CP-element group 136: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Update/ca
      -- 
    ca_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1033_inst_ack_1, ack => convolution3D_CP_1115_elements(136)); -- 
    -- CP-element group 137:  branch  join  transition  place  output  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	134 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (10) 
      -- CP-element group 137: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039__exit__
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040__entry__
      -- CP-element group 137: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/$exit
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_dead_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_eval_test/$entry
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_eval_test/$exit
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_eval_test/branch_req
      -- CP-element group 137: 	 branch_block_stmt_441/R_cmpx_xi_1041_place
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_if_link/$entry
      -- CP-element group 137: 	 branch_block_stmt_441/if_stmt_1040_else_link/$entry
      -- 
    branch_req_2214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(137), ack => if_stmt_1040_branch_req_0); -- 
    convolution3D_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(134) & convolution3D_CP_1115_elements(136);
      gj_convolution3D_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  place  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	320 
    -- CP-element group 138: 	321 
    -- CP-element group 138: 	323 
    -- CP-element group 138: 	324 
    -- CP-element group 138:  members (20) 
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/if_stmt_1040_if_link/$exit
      -- CP-element group 138: 	 branch_block_stmt_441/if_stmt_1040_if_link/if_choice_transition
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Update/cr
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Sample/rr
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Sample/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/$entry
      -- CP-element group 138: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/$entry
      -- 
    if_choice_transition_2219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1040_branch_ack_1, ack => convolution3D_CP_1115_elements(138)); -- 
    rr_3648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(138), ack => type_cast_992_inst_req_0); -- 
    cr_3653_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3653_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(138), ack => type_cast_992_inst_req_1); -- 
    cr_3676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(138), ack => type_cast_999_inst_req_1); -- 
    rr_3671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(138), ack => type_cast_999_inst_req_0); -- 
    -- CP-element group 139:  fork  transition  place  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	331 
    -- CP-element group 139: 	332 
    -- CP-element group 139:  members (12) 
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/if_stmt_1040_else_link/$exit
      -- CP-element group 139: 	 branch_block_stmt_441/if_stmt_1040_else_link/else_choice_transition
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Update/$entry
      -- CP-element group 139: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1040_branch_ack_0, ack => convolution3D_CP_1115_elements(139)); -- 
    rr_3707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(139), ack => type_cast_1050_inst_req_0); -- 
    cr_3712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(139), ack => type_cast_1050_inst_req_1); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	334 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	146 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_sample_complete
      -- CP-element group 140: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Sample/ack
      -- 
    ack_2254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_0, ack => convolution3D_CP_1115_elements(140)); -- 
    -- CP-element group 141:  transition  input  output  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	334 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	142 
    -- CP-element group 141:  members (11) 
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_offset_calculated
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Update/ack
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_request/$entry
      -- CP-element group 141: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_request/req
      -- 
    ack_2259_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1079_index_offset_ack_1, ack => convolution3D_CP_1115_elements(141)); -- 
    req_2268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(141), ack => addr_of_1080_final_reg_req_0); -- 
    -- CP-element group 142:  transition  input  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	141 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_request/$exit
      -- CP-element group 142: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_request/ack
      -- 
    ack_2269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_0, ack => convolution3D_CP_1115_elements(142)); -- 
    -- CP-element group 143:  join  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	334 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143:  members (28) 
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_complete/$exit
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_complete/ack
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_word_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_root_address_calculated
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_address_resized
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_addr_resize/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_addr_resize/$exit
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_addr_resize/base_resize_req
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_addr_resize/base_resize_ack
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_plus_offset/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_plus_offset/$exit
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_plus_offset/sum_rename_req
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_base_plus_offset/sum_rename_ack
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_word_addrgen/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_word_addrgen/$exit
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_word_addrgen/root_register_req
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_word_addrgen/root_register_ack
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/ptr_deref_1083_Split/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/ptr_deref_1083_Split/$exit
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/ptr_deref_1083_Split/split_req
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/ptr_deref_1083_Split/split_ack
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/word_0/rr
      -- 
    ack_2274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1080_final_reg_ack_1, ack => convolution3D_CP_1115_elements(143)); -- 
    rr_2312_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2312_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(143), ack => ptr_deref_1083_store_0_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/word_0/$exit
      -- CP-element group 144: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Sample/word_access_start/word_0/ra
      -- 
    ra_2313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1083_store_0_ack_0, ack => convolution3D_CP_1115_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	334 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	146 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/word_0/ca
      -- 
    ca_2324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1083_store_0_ack_1, ack => convolution3D_CP_1115_elements(145)); -- 
    -- CP-element group 146:  join  transition  place  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	140 
    -- CP-element group 146: 	145 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	335 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085__exit__
      -- CP-element group 146: 	 branch_block_stmt_441/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 146: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/$exit
      -- CP-element group 146: 	 branch_block_stmt_441/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- CP-element group 146: 	 branch_block_stmt_441/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(140) & convolution3D_CP_1115_elements(145);
      gj_convolution3D_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	335 
    -- CP-element group 147: successors 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Sample/ra
      -- 
    ra_2336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_0, ack => convolution3D_CP_1115_elements(147)); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	335 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	155 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Update/ca
      -- 
    ca_2341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1090_inst_ack_1, ack => convolution3D_CP_1115_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	335 
    -- CP-element group 149: successors 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Sample/ra
      -- 
    ra_2350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1094_inst_ack_0, ack => convolution3D_CP_1115_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	335 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	155 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Update/ca
      -- 
    ca_2355_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1094_inst_ack_1, ack => convolution3D_CP_1115_elements(150)); -- 
    -- CP-element group 151:  transition  input  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	335 
    -- CP-element group 151: successors 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Sample/ra
      -- 
    ra_2364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_0, ack => convolution3D_CP_1115_elements(151)); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	335 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	155 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Update/ca
      -- 
    ca_2369_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1098_inst_ack_1, ack => convolution3D_CP_1115_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	335 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Sample/ra
      -- 
    ra_2378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_0, ack => convolution3D_CP_1115_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	335 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Update/ca
      -- 
    ca_2383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1102_inst_ack_1, ack => convolution3D_CP_1115_elements(154)); -- 
    -- CP-element group 155:  branch  join  transition  place  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	148 
    -- CP-element group 155: 	150 
    -- CP-element group 155: 	152 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (10) 
      -- CP-element group 155: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139__exit__
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140__entry__
      -- CP-element group 155: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/$exit
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_dead_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_eval_test/$entry
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_eval_test/$exit
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_eval_test/branch_req
      -- CP-element group 155: 	 branch_block_stmt_441/R_cmp161379_1141_place
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_if_link/$entry
      -- CP-element group 155: 	 branch_block_stmt_441/if_stmt_1140_else_link/$entry
      -- 
    branch_req_2391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(155), ack => if_stmt_1140_branch_req_0); -- 
    convolution3D_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(148) & convolution3D_CP_1115_elements(150) & convolution3D_CP_1115_elements(152) & convolution3D_CP_1115_elements(154);
      gj_convolution3D_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156: 	159 
    -- CP-element group 156: 	160 
    -- CP-element group 156: 	161 
    -- CP-element group 156: 	162 
    -- CP-element group 156: 	163 
    -- CP-element group 156: 	164 
    -- CP-element group 156: 	165 
    -- CP-element group 156: 	168 
    -- CP-element group 156: 	170 
    -- CP-element group 156:  members (42) 
      -- CP-element group 156: 	 branch_block_stmt_441/merge_stmt_1146__exit__
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217__entry__
      -- CP-element group 156: 	 branch_block_stmt_441/merge_stmt_1146_PhiReqMerge
      -- CP-element group 156: 	 branch_block_stmt_441/if_stmt_1140_if_link/$exit
      -- CP-element group 156: 	 branch_block_stmt_441/if_stmt_1140_if_link/if_choice_transition
      -- CP-element group 156: 	 branch_block_stmt_441/ifx_xend_bbx_xnph
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_sample_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Sample/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Sample/rr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_update_start_
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Update/cr
      -- CP-element group 156: 	 branch_block_stmt_441/ifx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/ifx_xend_bbx_xnph_PhiReq/$exit
      -- CP-element group 156: 	 branch_block_stmt_441/merge_stmt_1146_PhiAck/$entry
      -- CP-element group 156: 	 branch_block_stmt_441/merge_stmt_1146_PhiAck/$exit
      -- CP-element group 156: 	 branch_block_stmt_441/merge_stmt_1146_PhiAck/dummy
      -- 
    if_choice_transition_2396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1140_branch_ack_1, ack => convolution3D_CP_1115_elements(156)); -- 
    rr_2413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1161_inst_req_0); -- 
    cr_2418_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2418_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1161_inst_req_1); -- 
    rr_2427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1165_inst_req_0); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1165_inst_req_1); -- 
    rr_2441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1174_inst_req_0); -- 
    cr_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1174_inst_req_1); -- 
    rr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1183_inst_req_0); -- 
    cr_2460_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2460_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1183_inst_req_1); -- 
    cr_2474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1192_inst_req_1); -- 
    cr_2488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(156), ack => type_cast_1197_inst_req_1); -- 
    -- CP-element group 157:  transition  place  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	345 
    -- CP-element group 157:  members (6) 
      -- CP-element group 157: 	 branch_block_stmt_441/if_stmt_1140_else_link/$exit
      -- CP-element group 157: 	 branch_block_stmt_441/if_stmt_1140_else_link/else_choice_transition
      -- CP-element group 157: 	 branch_block_stmt_441/ifx_xend_forx_xend215
      -- CP-element group 157: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/$entry
      -- CP-element group 157: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/$entry
      -- CP-element group 157: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/$entry
      -- 
    else_choice_transition_2400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1140_branch_ack_0, ack => convolution3D_CP_1115_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Sample/ra
      -- 
    ra_2414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_0, ack => convolution3D_CP_1115_elements(158)); -- 
    -- CP-element group 159:  transition  input  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	156 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	166 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1161_Update/ca
      -- 
    ca_2419_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1161_inst_ack_1, ack => convolution3D_CP_1115_elements(159)); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	156 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Sample/ra
      -- 
    ra_2428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1165_inst_ack_0, ack => convolution3D_CP_1115_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	156 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	166 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1165_Update/ca
      -- 
    ca_2433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1165_inst_ack_1, ack => convolution3D_CP_1115_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	156 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Sample/ra
      -- 
    ra_2442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_0, ack => convolution3D_CP_1115_elements(162)); -- 
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	156 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1174_Update/ca
      -- 
    ca_2447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1174_inst_ack_1, ack => convolution3D_CP_1115_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	156 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Sample/ra
      -- 
    ra_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1183_inst_ack_0, ack => convolution3D_CP_1115_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	156 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1183_Update/ca
      -- 
    ca_2461_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1183_inst_ack_1, ack => convolution3D_CP_1115_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	159 
    -- CP-element group 166: 	161 
    -- CP-element group 166: 	163 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Sample/rr
      -- 
    rr_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(166), ack => type_cast_1192_inst_req_0); -- 
    convolution3D_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(159) & convolution3D_CP_1115_elements(161) & convolution3D_CP_1115_elements(163) & convolution3D_CP_1115_elements(165);
      gj_convolution3D_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Sample/ra
      -- 
    ra_2470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_0, ack => convolution3D_CP_1115_elements(167)); -- 
    -- CP-element group 168:  transition  input  output  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	156 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	169 
    -- CP-element group 168:  members (6) 
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1192_Update/ca
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_sample_start_
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Sample/$entry
      -- CP-element group 168: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Sample/rr
      -- 
    ca_2475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1192_inst_ack_1, ack => convolution3D_CP_1115_elements(168)); -- 
    rr_2483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(168), ack => type_cast_1197_inst_req_0); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	168 
    -- CP-element group 169: successors 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Sample/ra
      -- 
    ra_2484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_0, ack => convolution3D_CP_1115_elements(169)); -- 
    -- CP-element group 170:  transition  place  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	156 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	336 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217__exit__
      -- CP-element group 170: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163
      -- CP-element group 170: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/$exit
      -- CP-element group 170: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_441/assign_stmt_1152_to_assign_stmt_1217/type_cast_1197_Update/ca
      -- CP-element group 170: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/$entry
      -- CP-element group 170: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/$entry
      -- CP-element group 170: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/$entry
      -- 
    ca_2489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_1, ack => convolution3D_CP_1115_elements(170)); -- 
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	341 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	210 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_sample_complete
      -- CP-element group 171: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Sample/ack
      -- 
    ack_2518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1232_index_offset_ack_0, ack => convolution3D_CP_1115_elements(171)); -- 
    -- CP-element group 172:  transition  input  output  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	341 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (11) 
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_root_address_calculated
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_offset_calculated
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_request/req
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_request/$entry
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_base_plus_offset/sum_rename_ack
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_base_plus_offset/sum_rename_req
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_base_plus_offset/$exit
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_base_plus_offset/$entry
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Update/ack
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_sample_start_
      -- 
    ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1232_index_offset_ack_1, ack => convolution3D_CP_1115_elements(172)); -- 
    req_2532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(172), ack => addr_of_1233_final_reg_req_0); -- 
    -- CP-element group 173:  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_request/ack
      -- CP-element group 173: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_request/$exit
      -- CP-element group 173: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_sample_completed_
      -- 
    ack_2533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1233_final_reg_ack_0, ack => convolution3D_CP_1115_elements(173)); -- 
    -- CP-element group 174:  fork  transition  input  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	341 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	207 
    -- CP-element group 174:  members (19) 
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_complete/ack
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_complete/$exit
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_word_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_root_address_calculated
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_address_resized
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_addr_resize/$entry
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_addr_resize/$exit
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_addr_resize/base_resize_req
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_addr_resize/base_resize_ack
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_plus_offset/$entry
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_plus_offset/$exit
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_plus_offset/sum_rename_req
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_base_plus_offset/sum_rename_ack
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_word_addrgen/$entry
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_word_addrgen/$exit
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_word_addrgen/root_register_req
      -- CP-element group 174: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_word_addrgen/root_register_ack
      -- 
    ack_2538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1233_final_reg_ack_1, ack => convolution3D_CP_1115_elements(174)); -- 
    -- CP-element group 175:  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	341 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175:  members (6) 
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Update/cr
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_update_start_
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Sample/ra
      -- CP-element group 175: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Update/$entry
      -- 
    ra_2547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1236_inst_ack_0, ack => convolution3D_CP_1115_elements(175)); -- 
    cr_2551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(175), ack => RPIPE_maxpool_input_pipe_1236_inst_req_1); -- 
    -- CP-element group 176:  fork  transition  input  output  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	177 
    -- CP-element group 176: 	179 
    -- CP-element group 176:  members (9) 
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Update/ca
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Sample/$entry
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_sample_start_
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Sample/rr
      -- CP-element group 176: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Sample/$entry
      -- 
    ca_2552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1236_inst_ack_1, ack => convolution3D_CP_1115_elements(176)); -- 
    rr_2560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(176), ack => type_cast_1240_inst_req_0); -- 
    rr_2574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(176), ack => RPIPE_maxpool_input_pipe_1249_inst_req_0); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	176 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_sample_completed_
      -- CP-element group 177: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Sample/ra
      -- CP-element group 177: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Sample/$exit
      -- 
    ra_2561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_0, ack => convolution3D_CP_1115_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	341 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	207 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Update/ca
      -- CP-element group 178: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Update/$exit
      -- 
    ca_2566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1240_inst_ack_1, ack => convolution3D_CP_1115_elements(178)); -- 
    -- CP-element group 179:  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	176 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179:  members (6) 
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Sample/ra
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_update_start_
      -- CP-element group 179: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_sample_completed_
      -- 
    ra_2575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1249_inst_ack_0, ack => convolution3D_CP_1115_elements(179)); -- 
    cr_2579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(179), ack => RPIPE_maxpool_input_pipe_1249_inst_req_1); -- 
    -- CP-element group 180:  fork  transition  input  output  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	181 
    -- CP-element group 180: 	183 
    -- CP-element group 180:  members (9) 
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Sample/rr
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Sample/$entry
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_sample_start_
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Update/ca
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1249_update_completed_
      -- 
    ca_2580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1249_inst_ack_1, ack => convolution3D_CP_1115_elements(180)); -- 
    rr_2588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(180), ack => type_cast_1253_inst_req_0); -- 
    rr_2602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(180), ack => RPIPE_maxpool_input_pipe_1267_inst_req_0); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	180 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Sample/ra
      -- CP-element group 181: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_sample_completed_
      -- 
    ra_2589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_0, ack => convolution3D_CP_1115_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	341 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	207 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Update/ca
      -- CP-element group 182: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Update/$exit
      -- CP-element group 182: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_update_completed_
      -- 
    ca_2594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1253_inst_ack_1, ack => convolution3D_CP_1115_elements(182)); -- 
    -- CP-element group 183:  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	180 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183:  members (6) 
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Update/cr
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_update_start_
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Sample/ra
      -- CP-element group 183: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Update/$entry
      -- 
    ra_2603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1267_inst_ack_0, ack => convolution3D_CP_1115_elements(183)); -- 
    cr_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(183), ack => RPIPE_maxpool_input_pipe_1267_inst_req_1); -- 
    -- CP-element group 184:  fork  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184: 	187 
    -- CP-element group 184:  members (9) 
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Update/ca
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1267_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Sample/rr
      -- CP-element group 184: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Sample/$entry
      -- 
    ca_2608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1267_inst_ack_1, ack => convolution3D_CP_1115_elements(184)); -- 
    rr_2616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(184), ack => type_cast_1271_inst_req_0); -- 
    rr_2630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(184), ack => RPIPE_maxpool_input_pipe_1285_inst_req_0); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Sample/$exit
      -- 
    ra_2617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_0, ack => convolution3D_CP_1115_elements(185)); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	341 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	207 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Update/ca
      -- CP-element group 186: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_update_completed_
      -- 
    ca_2622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1271_inst_ack_1, ack => convolution3D_CP_1115_elements(186)); -- 
    -- CP-element group 187:  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	184 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187:  members (6) 
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Update/cr
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Sample/ra
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_update_start_
      -- CP-element group 187: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_sample_completed_
      -- 
    ra_2631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1285_inst_ack_0, ack => convolution3D_CP_1115_elements(187)); -- 
    cr_2635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(187), ack => RPIPE_maxpool_input_pipe_1285_inst_req_1); -- 
    -- CP-element group 188:  fork  transition  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	189 
    -- CP-element group 188: 	191 
    -- CP-element group 188:  members (9) 
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_sample_start_
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Update/ca
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1285_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_sample_start_
      -- 
    ca_2636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1285_inst_ack_1, ack => convolution3D_CP_1115_elements(188)); -- 
    rr_2644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(188), ack => type_cast_1289_inst_req_0); -- 
    rr_2658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(188), ack => RPIPE_maxpool_input_pipe_1303_inst_req_0); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	188 
    -- CP-element group 189: successors 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Sample/ra
      -- 
    ra_2645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_0, ack => convolution3D_CP_1115_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	341 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	207 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Update/ca
      -- CP-element group 190: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Update/$exit
      -- 
    ca_2650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_1, ack => convolution3D_CP_1115_elements(190)); -- 
    -- CP-element group 191:  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	188 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191:  members (6) 
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Update/cr
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Sample/ra
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_update_start_
      -- CP-element group 191: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_sample_completed_
      -- 
    ra_2659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1303_inst_ack_0, ack => convolution3D_CP_1115_elements(191)); -- 
    cr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(191), ack => RPIPE_maxpool_input_pipe_1303_inst_req_1); -- 
    -- CP-element group 192:  fork  transition  input  output  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: 	195 
    -- CP-element group 192:  members (9) 
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Sample/$entry
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_Update/ca
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_sample_start_
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1303_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Sample/rr
      -- CP-element group 192: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Sample/$entry
      -- 
    ca_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1303_inst_ack_1, ack => convolution3D_CP_1115_elements(192)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(192), ack => type_cast_1307_inst_req_0); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(192), ack => RPIPE_maxpool_input_pipe_1321_inst_req_0); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	192 
    -- CP-element group 193: successors 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Sample/ra
      -- CP-element group 193: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_sample_completed_
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1307_inst_ack_0, ack => convolution3D_CP_1115_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	341 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	207 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Update/ca
      -- CP-element group 194: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_update_completed_
      -- 
    ca_2678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1307_inst_ack_1, ack => convolution3D_CP_1115_elements(194)); -- 
    -- CP-element group 195:  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	192 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (6) 
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Sample/$exit
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_sample_completed_
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Sample/ra
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_update_start_
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Update/cr
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1321_inst_ack_0, ack => convolution3D_CP_1115_elements(195)); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(195), ack => RPIPE_maxpool_input_pipe_1321_inst_req_1); -- 
    -- CP-element group 196:  fork  transition  input  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: 	199 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_update_completed_
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Sample/rr
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Update/ca
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1321_Update/$exit
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1321_inst_ack_1, ack => convolution3D_CP_1115_elements(196)); -- 
    rr_2700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(196), ack => type_cast_1325_inst_req_0); -- 
    rr_2714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(196), ack => RPIPE_maxpool_input_pipe_1339_inst_req_0); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Sample/ra
      -- CP-element group 197: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_sample_completed_
      -- 
    ra_2701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_0, ack => convolution3D_CP_1115_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	341 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	207 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Update/ca
      -- CP-element group 198: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_update_completed_
      -- 
    ca_2706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1325_inst_ack_1, ack => convolution3D_CP_1115_elements(198)); -- 
    -- CP-element group 199:  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	196 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199:  members (6) 
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Update/cr
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Sample/ra
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Sample/$exit
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_update_start_
      -- CP-element group 199: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_sample_completed_
      -- 
    ra_2715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1339_inst_ack_0, ack => convolution3D_CP_1115_elements(199)); -- 
    cr_2719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(199), ack => RPIPE_maxpool_input_pipe_1339_inst_req_1); -- 
    -- CP-element group 200:  fork  transition  input  output  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200: 	203 
    -- CP-element group 200:  members (9) 
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Update/ca
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_Update/$exit
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1339_update_completed_
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Sample/rr
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Sample/rr
      -- 
    ca_2720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1339_inst_ack_1, ack => convolution3D_CP_1115_elements(200)); -- 
    rr_2728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(200), ack => type_cast_1343_inst_req_0); -- 
    rr_2742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(200), ack => RPIPE_maxpool_input_pipe_1357_inst_req_0); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Sample/ra
      -- CP-element group 201: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_sample_completed_
      -- 
    ra_2729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_0, ack => convolution3D_CP_1115_elements(201)); -- 
    -- CP-element group 202:  transition  input  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	341 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	207 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Update/ca
      -- CP-element group 202: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_update_completed_
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1343_inst_ack_1, ack => convolution3D_CP_1115_elements(202)); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	200 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_update_start_
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_sample_completed_
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Sample/$exit
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Sample/ra
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Update/cr
      -- 
    ra_2743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1357_inst_ack_0, ack => convolution3D_CP_1115_elements(203)); -- 
    cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(203), ack => RPIPE_maxpool_input_pipe_1357_inst_req_1); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_update_completed_
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Update/$exit
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1357_Update/ca
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_sample_start_
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Sample/$entry
      -- CP-element group 204: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Sample/rr
      -- 
    ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1357_inst_ack_1, ack => convolution3D_CP_1115_elements(204)); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(204), ack => type_cast_1361_inst_req_0); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Sample/ra
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_0, ack => convolution3D_CP_1115_elements(205)); -- 
    -- CP-element group 206:  transition  input  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	341 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Update/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1361_inst_ack_1, ack => convolution3D_CP_1115_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	174 
    -- CP-element group 207: 	178 
    -- CP-element group 207: 	182 
    -- CP-element group 207: 	186 
    -- CP-element group 207: 	190 
    -- CP-element group 207: 	194 
    -- CP-element group 207: 	198 
    -- CP-element group 207: 	202 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (9) 
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/ptr_deref_1369_Split/$entry
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/ptr_deref_1369_Split/$exit
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/ptr_deref_1369_Split/split_req
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/ptr_deref_1369_Split/split_ack
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/$entry
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/word_0/$entry
      -- CP-element group 207: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/word_0/rr
      -- 
    rr_2800_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2800_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(207), ack => ptr_deref_1369_store_0_req_0); -- 
    convolution3D_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(174) & convolution3D_CP_1115_elements(178) & convolution3D_CP_1115_elements(182) & convolution3D_CP_1115_elements(186) & convolution3D_CP_1115_elements(190) & convolution3D_CP_1115_elements(194) & convolution3D_CP_1115_elements(198) & convolution3D_CP_1115_elements(202) & convolution3D_CP_1115_elements(206);
      gj_convolution3D_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/$exit
      -- CP-element group 208: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Sample/word_access_start/word_0/ra
      -- 
    ra_2801_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1369_store_0_ack_0, ack => convolution3D_CP_1115_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	341 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209:  members (5) 
      -- CP-element group 209: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/$exit
      -- CP-element group 209: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/word_0/$exit
      -- CP-element group 209: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/word_0/ca
      -- 
    ca_2812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1369_store_0_ack_1, ack => convolution3D_CP_1115_elements(209)); -- 
    -- CP-element group 210:  branch  join  transition  place  output  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	171 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	211 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (10) 
      -- CP-element group 210: 	 branch_block_stmt_441/R_exitcond_1384_place
      -- CP-element group 210: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382__exit__
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383__entry__
      -- CP-element group 210: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/$exit
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_dead_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_eval_test/$entry
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_eval_test/$exit
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_eval_test/branch_req
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_if_link/$entry
      -- CP-element group 210: 	 branch_block_stmt_441/if_stmt_1383_else_link/$entry
      -- 
    branch_req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(210), ack => if_stmt_1383_branch_req_0); -- 
    convolution3D_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(171) & convolution3D_CP_1115_elements(209);
      gj_convolution3D_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	210 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	342 
    -- CP-element group 211: 	343 
    -- CP-element group 211:  members (24) 
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge
      -- CP-element group 211: 	 branch_block_stmt_441/merge_stmt_1389__exit__
      -- CP-element group 211: 	 branch_block_stmt_441/assign_stmt_1396_to_assign_stmt_1411__entry__
      -- CP-element group 211: 	 branch_block_stmt_441/assign_stmt_1396_to_assign_stmt_1411__exit__
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215
      -- CP-element group 211: 	 branch_block_stmt_441/merge_stmt_1389_PhiReqMerge
      -- CP-element group 211: 	 branch_block_stmt_441/if_stmt_1383_if_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_441/if_stmt_1383_if_link/if_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_441/assign_stmt_1396_to_assign_stmt_1411/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/assign_stmt_1396_to_assign_stmt_1411/$exit
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xbody163_forx_xcond156x_xforx_xend215_crit_edge_PhiReq/$exit
      -- CP-element group 211: 	 branch_block_stmt_441/merge_stmt_1389_PhiAck/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/merge_stmt_1389_PhiAck/$exit
      -- CP-element group 211: 	 branch_block_stmt_441/merge_stmt_1389_PhiAck/dummy
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_1, ack => convolution3D_CP_1115_elements(211)); -- 
    rr_3815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(211), ack => type_cast_1417_inst_req_0); -- 
    cr_3820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(211), ack => type_cast_1417_inst_req_1); -- 
    -- CP-element group 212:  fork  transition  place  input  output  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	337 
    -- CP-element group 212: 	338 
    -- CP-element group 212:  members (12) 
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163
      -- CP-element group 212: 	 branch_block_stmt_441/if_stmt_1383_else_link/$exit
      -- CP-element group 212: 	 branch_block_stmt_441/if_stmt_1383_else_link/else_choice_transition
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Sample/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Sample/rr
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1383_branch_ack_0, ack => convolution3D_CP_1115_elements(212)); -- 
    rr_3772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(212), ack => type_cast_1226_inst_req_0); -- 
    cr_3777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(212), ack => type_cast_1226_inst_req_1); -- 
    -- CP-element group 213:  transition  place  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	347 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	366 
    -- CP-element group 213:  members (5) 
      -- CP-element group 213: 	 branch_block_stmt_441/forx_xend215_ifx_xend227
      -- CP-element group 213: 	 branch_block_stmt_441/if_stmt_1434_if_link/$exit
      -- CP-element group 213: 	 branch_block_stmt_441/if_stmt_1434_if_link/if_choice_transition
      -- CP-element group 213: 	 branch_block_stmt_441/forx_xend215_ifx_xend227_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_441/forx_xend215_ifx_xend227_PhiReq/$exit
      -- 
    if_choice_transition_2850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1434_branch_ack_1, ack => convolution3D_CP_1115_elements(213)); -- 
    -- CP-element group 214:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	347 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (18) 
      -- CP-element group 214: 	 branch_block_stmt_441/forx_xend215_bbx_xnphx_xi356
      -- CP-element group 214: 	 branch_block_stmt_441/merge_stmt_1440__exit__
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456__entry__
      -- CP-element group 214: 	 branch_block_stmt_441/merge_stmt_1440_PhiReqMerge
      -- CP-element group 214: 	 branch_block_stmt_441/if_stmt_1434_else_link/$exit
      -- CP-element group 214: 	 branch_block_stmt_441/if_stmt_1434_else_link/else_choice_transition
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/$entry
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_update_start_
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Sample/rr
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Update/cr
      -- CP-element group 214: 	 branch_block_stmt_441/forx_xend215_bbx_xnphx_xi356_PhiReq/$entry
      -- CP-element group 214: 	 branch_block_stmt_441/forx_xend215_bbx_xnphx_xi356_PhiReq/$exit
      -- CP-element group 214: 	 branch_block_stmt_441/merge_stmt_1440_PhiAck/$entry
      -- CP-element group 214: 	 branch_block_stmt_441/merge_stmt_1440_PhiAck/$exit
      -- CP-element group 214: 	 branch_block_stmt_441/merge_stmt_1440_PhiAck/dummy
      -- 
    else_choice_transition_2854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1434_branch_ack_0, ack => convolution3D_CP_1115_elements(214)); -- 
    rr_2867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(214), ack => type_cast_1449_inst_req_0); -- 
    cr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(214), ack => type_cast_1449_inst_req_1); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Sample/ra
      -- 
    ra_2868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_0, ack => convolution3D_CP_1115_elements(215)); -- 
    -- CP-element group 216:  fork  transition  place  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	348 
    -- CP-element group 216: 	349 
    -- CP-element group 216:  members (11) 
      -- CP-element group 216: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456__exit__
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365
      -- CP-element group 216: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/$exit
      -- CP-element group 216: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_441/assign_stmt_1446_to_assign_stmt_1456/type_cast_1449_Update/ca
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/$entry
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/$entry
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/$entry
      -- CP-element group 216: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$entry
      -- 
    ca_2873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1449_inst_ack_1, ack => convolution3D_CP_1115_elements(216)); -- 
    -- CP-element group 217:  transition  input  output  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	361 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (6) 
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_sample_completed_
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_update_start_
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Sample/$exit
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Sample/ra
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Update/$entry
      -- CP-element group 217: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Update/cr
      -- 
    ra_2885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1487_inst_ack_0, ack => convolution3D_CP_1115_elements(217)); -- 
    cr_2889_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2889_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(217), ack => RPIPE_maxpool_input_pipe_1487_inst_req_1); -- 
    -- CP-element group 218:  transition  input  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218:  members (6) 
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_update_completed_
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Update/$exit
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Update/ca
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Sample/rr
      -- 
    ca_2890_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1487_inst_ack_1, ack => convolution3D_CP_1115_elements(218)); -- 
    rr_2898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(218), ack => type_cast_1491_inst_req_0); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Sample/ra
      -- 
    ra_2899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1491_inst_ack_0, ack => convolution3D_CP_1115_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	361 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	223 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Update/ca
      -- 
    ca_2904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1491_inst_ack_1, ack => convolution3D_CP_1115_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	361 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Sample/$exit
      -- CP-element group 221: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Sample/ra
      -- 
    ra_2913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1506_inst_ack_0, ack => convolution3D_CP_1115_elements(221)); -- 
    -- CP-element group 222:  transition  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	361 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Update/ca
      -- 
    ca_2918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1506_inst_ack_1, ack => convolution3D_CP_1115_elements(222)); -- 
    -- CP-element group 223:  branch  join  transition  place  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	220 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	224 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (10) 
      -- CP-element group 223: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512__exit__
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513__entry__
      -- CP-element group 223: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/$exit
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_dead_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_eval_test/$entry
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_eval_test/$exit
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_eval_test/branch_req
      -- CP-element group 223: 	 branch_block_stmt_441/R_cmpx_xi364_1514_place
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_if_link/$entry
      -- CP-element group 223: 	 branch_block_stmt_441/if_stmt_1513_else_link/$entry
      -- 
    branch_req_2926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(223), ack => if_stmt_1513_branch_req_0); -- 
    convolution3D_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(220) & convolution3D_CP_1115_elements(222);
      gj_convolution3D_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	223 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	351 
    -- CP-element group 224: 	352 
    -- CP-element group 224: 	354 
    -- CP-element group 224: 	355 
    -- CP-element group 224:  members (20) 
      -- CP-element group 224: 	 branch_block_stmt_441/if_stmt_1513_if_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_441/if_stmt_1513_if_link/if_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Update/cr
      -- 
    if_choice_transition_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1513_branch_ack_1, ack => convolution3D_CP_1115_elements(224)); -- 
    rr_3888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(224), ack => type_cast_1465_inst_req_0); -- 
    cr_3893_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3893_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(224), ack => type_cast_1465_inst_req_1); -- 
    rr_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(224), ack => type_cast_1472_inst_req_0); -- 
    cr_3916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(224), ack => type_cast_1472_inst_req_1); -- 
    -- CP-element group 225:  fork  transition  place  input  output  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	362 
    -- CP-element group 225: 	363 
    -- CP-element group 225:  members (12) 
      -- CP-element group 225: 	 branch_block_stmt_441/if_stmt_1513_else_link/$exit
      -- CP-element group 225: 	 branch_block_stmt_441/if_stmt_1513_else_link/else_choice_transition
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Sample/rr
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Update/$entry
      -- CP-element group 225: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1513_branch_ack_0, ack => convolution3D_CP_1115_elements(225)); -- 
    rr_3947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(225), ack => type_cast_1523_inst_req_0); -- 
    cr_3952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(225), ack => type_cast_1523_inst_req_1); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	365 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	232 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_sample_complete
      -- CP-element group 226: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Sample/$exit
      -- CP-element group 226: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Sample/ack
      -- 
    ack_2966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1552_index_offset_ack_0, ack => convolution3D_CP_1115_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	365 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (11) 
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_sample_start_
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_root_address_calculated
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_offset_calculated
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Update/$exit
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Update/ack
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_base_plus_offset/$entry
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_base_plus_offset/$exit
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_base_plus_offset/sum_rename_req
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_base_plus_offset/sum_rename_ack
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_request/$entry
      -- CP-element group 227: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_request/req
      -- 
    ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1552_index_offset_ack_1, ack => convolution3D_CP_1115_elements(227)); -- 
    req_2980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(227), ack => addr_of_1553_final_reg_req_0); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_request/$exit
      -- CP-element group 228: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_request/ack
      -- 
    ack_2981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1553_final_reg_ack_0, ack => convolution3D_CP_1115_elements(228)); -- 
    -- CP-element group 229:  join  fork  transition  input  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	365 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (28) 
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_complete/$exit
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_complete/ack
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_word_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_root_address_calculated
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_address_resized
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_addr_resize/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_addr_resize/$exit
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_addr_resize/base_resize_req
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_addr_resize/base_resize_ack
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_plus_offset/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_plus_offset/$exit
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_plus_offset/sum_rename_req
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_base_plus_offset/sum_rename_ack
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_word_addrgen/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_word_addrgen/$exit
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_word_addrgen/root_register_req
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_word_addrgen/root_register_ack
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/ptr_deref_1556_Split/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/ptr_deref_1556_Split/$exit
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/ptr_deref_1556_Split/split_req
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/ptr_deref_1556_Split/split_ack
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/word_0/$entry
      -- CP-element group 229: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/word_0/rr
      -- 
    ack_2986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1553_final_reg_ack_1, ack => convolution3D_CP_1115_elements(229)); -- 
    rr_3024_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3024_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(229), ack => ptr_deref_1556_store_0_req_0); -- 
    -- CP-element group 230:  transition  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230:  members (5) 
      -- CP-element group 230: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/$exit
      -- CP-element group 230: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/word_0/$exit
      -- CP-element group 230: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Sample/word_access_start/word_0/ra
      -- 
    ra_3025_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1556_store_0_ack_0, ack => convolution3D_CP_1115_elements(230)); -- 
    -- CP-element group 231:  transition  input  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	365 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231:  members (5) 
      -- CP-element group 231: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/$exit
      -- CP-element group 231: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/word_0/$exit
      -- CP-element group 231: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/word_0/ca
      -- 
    ca_3036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1556_store_0_ack_1, ack => convolution3D_CP_1115_elements(231)); -- 
    -- CP-element group 232:  join  transition  place  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	226 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	366 
    -- CP-element group 232:  members (5) 
      -- CP-element group 232: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558__exit__
      -- CP-element group 232: 	 branch_block_stmt_441/getRemainingElementsx_xexit373_ifx_xend227
      -- CP-element group 232: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/$exit
      -- CP-element group 232: 	 branch_block_stmt_441/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$entry
      -- CP-element group 232: 	 branch_block_stmt_441/getRemainingElementsx_xexit373_ifx_xend227_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_232: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_232"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(226) & convolution3D_CP_1115_elements(231);
      gj_convolution3D_cp_element_group_232 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(232), clk => clk, reset => reset); --
    end block;
    -- CP-element group 233:  transition  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	366 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_sample_completed_
      -- CP-element group 233: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Sample/$exit
      -- CP-element group 233: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Sample/cra
      -- 
    cra_3048_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1563_call_ack_0, ack => convolution3D_CP_1115_elements(233)); -- 
    -- CP-element group 234:  fork  transition  place  input  output  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	366 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	235 
    -- CP-element group 234: 	237 
    -- CP-element group 234: 	241 
    -- CP-element group 234: 	242 
    -- CP-element group 234: 	243 
    -- CP-element group 234: 	244 
    -- CP-element group 234: 	245 
    -- CP-element group 234: 	246 
    -- CP-element group 234:  members (31) 
      -- CP-element group 234: 	 branch_block_stmt_441/call_stmt_1563__exit__
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631__entry__
      -- CP-element group 234: 	 branch_block_stmt_441/call_stmt_1563/$exit
      -- CP-element group 234: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_update_completed_
      -- CP-element group 234: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Update/$exit
      -- CP-element group 234: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Update/cca
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Sample/req
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_update_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_update_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Update/cr
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_update_start_
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Sample/rr
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Update/cr
      -- 
    cca_3053_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1563_call_ack_1, ack => convolution3D_CP_1115_elements(234)); -- 
    req_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => WPIPE_num_out_pipe_1575_inst_req_0); -- 
    req_3078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => WPIPE_maxpool_output_pipe_1578_inst_req_0); -- 
    rr_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1606_inst_req_0); -- 
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1606_inst_req_1); -- 
    rr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1616_inst_req_0); -- 
    cr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1616_inst_req_1); -- 
    rr_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1625_inst_req_0); -- 
    cr_3139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(234), ack => type_cast_1625_inst_req_1); -- 
    -- CP-element group 235:  transition  input  output  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	234 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (6) 
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_update_start_
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Sample/ack
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Update/req
      -- 
    ack_3065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1575_inst_ack_0, ack => convolution3D_CP_1115_elements(235)); -- 
    req_3069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(235), ack => WPIPE_num_out_pipe_1575_inst_req_1); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	247 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_num_out_pipe_1575_Update/ack
      -- 
    ack_3070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1575_inst_ack_1, ack => convolution3D_CP_1115_elements(236)); -- 
    -- CP-element group 237:  transition  input  output  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	234 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	238 
    -- CP-element group 237:  members (6) 
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_sample_completed_
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_update_start_
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Sample/ack
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Update/$entry
      -- CP-element group 237: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Update/req
      -- 
    ack_3079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1578_inst_ack_0, ack => convolution3D_CP_1115_elements(237)); -- 
    req_3083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(237), ack => WPIPE_maxpool_output_pipe_1578_inst_req_1); -- 
    -- CP-element group 238:  transition  input  output  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	237 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (6) 
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_update_completed_
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1578_Update/ack
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Sample/req
      -- 
    ack_3084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1578_inst_ack_1, ack => convolution3D_CP_1115_elements(238)); -- 
    req_3092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(238), ack => WPIPE_maxpool_output_pipe_1582_inst_req_0); -- 
    -- CP-element group 239:  transition  input  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (6) 
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_update_start_
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Sample/ack
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Update/req
      -- 
    ack_3093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_0, ack => convolution3D_CP_1115_elements(239)); -- 
    req_3097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(239), ack => WPIPE_maxpool_output_pipe_1582_inst_req_1); -- 
    -- CP-element group 240:  transition  input  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	247 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/WPIPE_maxpool_output_pipe_1582_Update/ack
      -- 
    ack_3098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1582_inst_ack_1, ack => convolution3D_CP_1115_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	234 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Sample/ra
      -- 
    ra_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_0, ack => convolution3D_CP_1115_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	234 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	247 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1606_Update/ca
      -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1606_inst_ack_1, ack => convolution3D_CP_1115_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	234 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Sample/ra
      -- 
    ra_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1616_inst_ack_0, ack => convolution3D_CP_1115_elements(243)); -- 
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	234 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	247 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1616_Update/ca
      -- 
    ca_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1616_inst_ack_1, ack => convolution3D_CP_1115_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	234 
    -- CP-element group 245: successors 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_sample_completed_
      -- CP-element group 245: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Sample/$exit
      -- CP-element group 245: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Sample/ra
      -- 
    ra_3135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_0, ack => convolution3D_CP_1115_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	234 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_update_completed_
      -- CP-element group 246: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Update/$exit
      -- CP-element group 246: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/type_cast_1625_Update/ca
      -- 
    ca_3140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1625_inst_ack_1, ack => convolution3D_CP_1115_elements(246)); -- 
    -- CP-element group 247:  join  transition  place  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	236 
    -- CP-element group 247: 	240 
    -- CP-element group 247: 	242 
    -- CP-element group 247: 	244 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	367 
    -- CP-element group 247:  members (6) 
      -- CP-element group 247: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631__exit__
      -- CP-element group 247: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody
      -- CP-element group 247: 	 branch_block_stmt_441/assign_stmt_1569_to_assign_stmt_1631/$exit
      -- CP-element group 247: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/$entry
      -- CP-element group 247: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/$entry
      -- CP-element group 247: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/$entry
      -- 
    convolution3D_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(236) & convolution3D_CP_1115_elements(240) & convolution3D_CP_1115_elements(242) & convolution3D_CP_1115_elements(244) & convolution3D_CP_1115_elements(246);
      gj_convolution3D_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	372 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Sample/ra
      -- 
    ra_3152_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1654_inst_ack_0, ack => convolution3D_CP_1115_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	372 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	252 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Update/ca
      -- 
    ca_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1654_inst_ack_1, ack => convolution3D_CP_1115_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	372 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Sample/ra
      -- 
    ra_3166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_0, ack => convolution3D_CP_1115_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	372 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Update/ca
      -- 
    ca_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1658_inst_ack_1, ack => convolution3D_CP_1115_elements(251)); -- 
    -- CP-element group 252:  join  transition  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	249 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_sample_start_
      -- CP-element group 252: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Sample/$entry
      -- CP-element group 252: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Sample/crr
      -- 
    crr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(252), ack => call_stmt_1662_call_req_0); -- 
    convolution3D_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(249) & convolution3D_CP_1115_elements(251);
      gj_convolution3D_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_sample_completed_
      -- CP-element group 253: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Sample/$exit
      -- CP-element group 253: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Sample/cra
      -- 
    cra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1662_call_ack_0, ack => convolution3D_CP_1115_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	372 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	257 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_update_completed_
      -- CP-element group 254: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Update/$exit
      -- CP-element group 254: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Update/cca
      -- 
    cca_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1662_call_ack_1, ack => convolution3D_CP_1115_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	372 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Sample/cra
      -- 
    cra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1669_call_ack_0, ack => convolution3D_CP_1115_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	372 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	257 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Update/cca
      -- 
    cca_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1669_call_ack_1, ack => convolution3D_CP_1115_elements(256)); -- 
    -- CP-element group 257:  branch  join  transition  place  output  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	254 
    -- CP-element group 257: 	256 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	258 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (10) 
      -- CP-element group 257: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680__exit__
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681__entry__
      -- CP-element group 257: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/$exit
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_dead_link/$entry
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_eval_test/$entry
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_eval_test/$exit
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_eval_test/branch_req
      -- CP-element group 257: 	 branch_block_stmt_441/R_exitcond5_1682_place
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_if_link/$entry
      -- CP-element group 257: 	 branch_block_stmt_441/if_stmt_1681_else_link/$entry
      -- 
    branch_req_3207_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3207_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(257), ack => if_stmt_1681_branch_req_0); -- 
    convolution3D_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(254) & convolution3D_CP_1115_elements(256);
      gj_convolution3D_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	257 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	261 
    -- CP-element group 258:  members (18) 
      -- CP-element group 258: 	 branch_block_stmt_441/merge_stmt_1687__exit__
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692__entry__
      -- CP-element group 258: 	 branch_block_stmt_441/if_stmt_1681_if_link/$exit
      -- CP-element group 258: 	 branch_block_stmt_441/if_stmt_1681_if_link/if_choice_transition
      -- CP-element group 258: 	 branch_block_stmt_441/whilex_xbody_whilex_xend
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/$entry
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_update_start_
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Sample/rr
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Update/cr
      -- CP-element group 258: 	 branch_block_stmt_441/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 258: 	 branch_block_stmt_441/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 258: 	 branch_block_stmt_441/merge_stmt_1687_PhiReqMerge
      -- CP-element group 258: 	 branch_block_stmt_441/merge_stmt_1687_PhiAck/$entry
      -- CP-element group 258: 	 branch_block_stmt_441/merge_stmt_1687_PhiAck/$exit
      -- CP-element group 258: 	 branch_block_stmt_441/merge_stmt_1687_PhiAck/dummy
      -- 
    if_choice_transition_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1681_branch_ack_1, ack => convolution3D_CP_1115_elements(258)); -- 
    rr_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(258), ack => type_cast_1691_inst_req_0); -- 
    cr_3234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(258), ack => type_cast_1691_inst_req_1); -- 
    -- CP-element group 259:  fork  transition  place  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	368 
    -- CP-element group 259: 	369 
    -- CP-element group 259:  members (12) 
      -- CP-element group 259: 	 branch_block_stmt_441/if_stmt_1681_else_link/$exit
      -- CP-element group 259: 	 branch_block_stmt_441/if_stmt_1681_else_link/else_choice_transition
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Sample/rr
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1681_branch_ack_0, ack => convolution3D_CP_1115_elements(259)); -- 
    rr_4000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(259), ack => type_cast_1637_inst_req_0); -- 
    cr_4005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(259), ack => type_cast_1637_inst_req_1); -- 
    -- CP-element group 260:  transition  input  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Sample/ra
      -- 
    ra_3230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1691_inst_ack_0, ack => convolution3D_CP_1115_elements(260)); -- 
    -- CP-element group 261:  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	258 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261: 	263 
    -- CP-element group 261: 	265 
    -- CP-element group 261: 	267 
    -- CP-element group 261: 	269 
    -- CP-element group 261: 	271 
    -- CP-element group 261: 	273 
    -- CP-element group 261: 	275 
    -- CP-element group 261: 	277 
    -- CP-element group 261: 	279 
    -- CP-element group 261: 	281 
    -- CP-element group 261:  members (40) 
      -- CP-element group 261: 	 branch_block_stmt_441/assign_stmt_1692__exit__
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803__entry__
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/assign_stmt_1692/$exit
      -- CP-element group 261: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_441/assign_stmt_1692/type_cast_1691_Update/ca
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Sample/crr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Update/ccr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_update_start_
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Update/cr
      -- CP-element group 261: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_update_start_
      -- 
    ca_3235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1691_inst_ack_1, ack => convolution3D_CP_1115_elements(261)); -- 
    cr_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1778_inst_req_1); -- 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1748_inst_req_1); -- 
    cr_3349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1758_inst_req_1); -- 
    cr_3363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1768_inst_req_1); -- 
    crr_3246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => call_stmt_1695_call_req_0); -- 
    ccr_3251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => call_stmt_1695_call_req_1); -- 
    cr_3265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1699_inst_req_1); -- 
    cr_3279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1708_inst_req_1); -- 
    cr_3293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1718_inst_req_1); -- 
    cr_3307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1728_inst_req_1); -- 
    cr_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(261), ack => type_cast_1738_inst_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_sample_completed_
      -- CP-element group 262: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Sample/cra
      -- 
    cra_3247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1695_call_ack_0, ack => convolution3D_CP_1115_elements(262)); -- 
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_update_completed_
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/call_stmt_1695_Update/cca
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_sample_start_
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Sample/$entry
      -- CP-element group 263: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Sample/rr
      -- 
    cca_3252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1695_call_ack_1, ack => convolution3D_CP_1115_elements(263)); -- 
    rr_3260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(263), ack => type_cast_1699_inst_req_0); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Sample/ra
      -- 
    ra_3261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1699_inst_ack_0, ack => convolution3D_CP_1115_elements(264)); -- 
    -- CP-element group 265:  fork  transition  input  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	261 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265: 	268 
    -- CP-element group 265: 	270 
    -- CP-element group 265: 	272 
    -- CP-element group 265: 	274 
    -- CP-element group 265: 	276 
    -- CP-element group 265: 	278 
    -- CP-element group 265: 	280 
    -- CP-element group 265:  members (27) 
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1699_Update/ca
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_sample_start_
      -- 
    ca_3266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1699_inst_ack_1, ack => convolution3D_CP_1115_elements(265)); -- 
    rr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1708_inst_req_0); -- 
    rr_3288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1718_inst_req_0); -- 
    rr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1728_inst_req_0); -- 
    rr_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1738_inst_req_0); -- 
    rr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1748_inst_req_0); -- 
    rr_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1758_inst_req_0); -- 
    rr_3358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1768_inst_req_0); -- 
    rr_3372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(265), ack => type_cast_1778_inst_req_0); -- 
    -- CP-element group 266:  transition  input  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Sample/ra
      -- 
    ra_3275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_0, ack => convolution3D_CP_1115_elements(266)); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	261 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	302 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_update_completed_
      -- CP-element group 267: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1708_Update/ca
      -- 
    ca_3280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1708_inst_ack_1, ack => convolution3D_CP_1115_elements(267)); -- 
    -- CP-element group 268:  transition  input  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	265 
    -- CP-element group 268: successors 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Sample/ra
      -- 
    ra_3289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_0, ack => convolution3D_CP_1115_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	261 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	299 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1718_Update/ca
      -- 
    ca_3294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1718_inst_ack_1, ack => convolution3D_CP_1115_elements(269)); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	265 
    -- CP-element group 270: successors 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_sample_completed_
      -- CP-element group 270: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Sample/ra
      -- 
    ra_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_0, ack => convolution3D_CP_1115_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	261 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	296 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_update_completed_
      -- CP-element group 271: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1728_Update/ca
      -- 
    ca_3308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1728_inst_ack_1, ack => convolution3D_CP_1115_elements(271)); -- 
    -- CP-element group 272:  transition  input  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	265 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Sample/ra
      -- 
    ra_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_0, ack => convolution3D_CP_1115_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	261 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	293 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1738_Update/ca
      -- 
    ca_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1738_inst_ack_1, ack => convolution3D_CP_1115_elements(273)); -- 
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	265 
    -- CP-element group 274: successors 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Sample/ra
      -- CP-element group 274: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_sample_completed_
      -- 
    ra_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_0, ack => convolution3D_CP_1115_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	261 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	290 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_Update/ca
      -- CP-element group 275: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1748_update_completed_
      -- 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_1, ack => convolution3D_CP_1115_elements(275)); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	265 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_sample_completed_
      -- CP-element group 276: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Sample/ra
      -- 
    ra_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1758_inst_ack_0, ack => convolution3D_CP_1115_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	261 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	287 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Update/ca
      -- CP-element group 277: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_update_completed_
      -- CP-element group 277: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1758_Update/$exit
      -- 
    ca_3350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1758_inst_ack_1, ack => convolution3D_CP_1115_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	265 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Sample/ra
      -- CP-element group 278: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Sample/$exit
      -- 
    ra_3359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_0, ack => convolution3D_CP_1115_elements(278)); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	261 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	284 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Update/ca
      -- CP-element group 279: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1768_update_completed_
      -- 
    ca_3364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1768_inst_ack_1, ack => convolution3D_CP_1115_elements(279)); -- 
    -- CP-element group 280:  transition  input  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	265 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Sample/ra
      -- CP-element group 280: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_sample_completed_
      -- 
    ra_3373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1778_inst_ack_0, ack => convolution3D_CP_1115_elements(280)); -- 
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	261 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_Update/ca
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_sample_start_
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Sample/req
      -- CP-element group 281: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/type_cast_1778_update_completed_
      -- 
    ca_3378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1778_inst_ack_1, ack => convolution3D_CP_1115_elements(281)); -- 
    req_3386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(281), ack => WPIPE_maxpool_output_pipe_1780_inst_req_0); -- 
    -- CP-element group 282:  transition  input  output  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	283 
    -- CP-element group 282:  members (6) 
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_sample_completed_
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_update_start_
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Sample/$exit
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Sample/ack
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Update/req
      -- CP-element group 282: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Update/$entry
      -- 
    ack_3387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1780_inst_ack_0, ack => convolution3D_CP_1115_elements(282)); -- 
    req_3391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(282), ack => WPIPE_maxpool_output_pipe_1780_inst_req_1); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	282 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_update_completed_
      -- CP-element group 283: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Update/ack
      -- CP-element group 283: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1780_Update/$exit
      -- 
    ack_3392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1780_inst_ack_1, ack => convolution3D_CP_1115_elements(283)); -- 
    -- CP-element group 284:  join  transition  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	279 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	285 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Sample/req
      -- 
    req_3400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(284), ack => WPIPE_maxpool_output_pipe_1783_inst_req_0); -- 
    convolution3D_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(279) & convolution3D_CP_1115_elements(283);
      gj_convolution3D_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  output  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	284 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (6) 
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_sample_completed_
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_update_start_
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Update/req
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Update/$entry
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Sample/ack
      -- CP-element group 285: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Sample/$exit
      -- 
    ack_3401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1783_inst_ack_0, ack => convolution3D_CP_1115_elements(285)); -- 
    req_3405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(285), ack => WPIPE_maxpool_output_pipe_1783_inst_req_1); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_update_completed_
      -- CP-element group 286: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Update/ack
      -- CP-element group 286: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1783_Update/$exit
      -- 
    ack_3406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1783_inst_ack_1, ack => convolution3D_CP_1115_elements(286)); -- 
    -- CP-element group 287:  join  transition  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	277 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Sample/req
      -- CP-element group 287: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Sample/$entry
      -- CP-element group 287: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_sample_start_
      -- 
    req_3414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(287), ack => WPIPE_maxpool_output_pipe_1786_inst_req_0); -- 
    convolution3D_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(277) & convolution3D_CP_1115_elements(286);
      gj_convolution3D_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  transition  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	289 
    -- CP-element group 288:  members (6) 
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Update/req
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_update_start_
      -- CP-element group 288: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_sample_completed_
      -- 
    ack_3415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1786_inst_ack_0, ack => convolution3D_CP_1115_elements(288)); -- 
    req_3419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(288), ack => WPIPE_maxpool_output_pipe_1786_inst_req_1); -- 
    -- CP-element group 289:  transition  input  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	288 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	290 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Update/ack
      -- CP-element group 289: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1786_update_completed_
      -- 
    ack_3420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1786_inst_ack_1, ack => convolution3D_CP_1115_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	275 
    -- CP-element group 290: 	289 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	291 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Sample/req
      -- CP-element group 290: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_sample_start_
      -- 
    req_3428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(290), ack => WPIPE_maxpool_output_pipe_1789_inst_req_0); -- 
    convolution3D_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(275) & convolution3D_CP_1115_elements(289);
      gj_convolution3D_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  transition  input  output  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	290 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	292 
    -- CP-element group 291:  members (6) 
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Update/req
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Sample/ack
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_update_start_
      -- CP-element group 291: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_sample_completed_
      -- 
    ack_3429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1789_inst_ack_0, ack => convolution3D_CP_1115_elements(291)); -- 
    req_3433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(291), ack => WPIPE_maxpool_output_pipe_1789_inst_req_1); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	291 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Update/ack
      -- CP-element group 292: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1789_update_completed_
      -- 
    ack_3434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1789_inst_ack_1, ack => convolution3D_CP_1115_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	273 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Sample/req
      -- CP-element group 293: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_sample_start_
      -- 
    req_3442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(293), ack => WPIPE_maxpool_output_pipe_1792_inst_req_0); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(273) & convolution3D_CP_1115_elements(292);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  transition  input  output  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (6) 
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Update/$entry
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Update/req
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Sample/ack
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Sample/$exit
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_update_start_
      -- CP-element group 294: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_sample_completed_
      -- 
    ack_3443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1792_inst_ack_0, ack => convolution3D_CP_1115_elements(294)); -- 
    req_3447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(294), ack => WPIPE_maxpool_output_pipe_1792_inst_req_1); -- 
    -- CP-element group 295:  transition  input  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	296 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Update/$exit
      -- CP-element group 295: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_Update/ack
      -- CP-element group 295: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1792_update_completed_
      -- 
    ack_3448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1792_inst_ack_1, ack => convolution3D_CP_1115_elements(295)); -- 
    -- CP-element group 296:  join  transition  output  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	271 
    -- CP-element group 296: 	295 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	297 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_sample_start_
      -- CP-element group 296: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Sample/$entry
      -- CP-element group 296: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Sample/req
      -- 
    req_3456_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3456_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(296), ack => WPIPE_maxpool_output_pipe_1795_inst_req_0); -- 
    convolution3D_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(271) & convolution3D_CP_1115_elements(295);
      gj_convolution3D_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  transition  input  output  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	296 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (6) 
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_sample_completed_
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_update_start_
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Sample/ack
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Update/$entry
      -- CP-element group 297: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Update/req
      -- 
    ack_3457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1795_inst_ack_0, ack => convolution3D_CP_1115_elements(297)); -- 
    req_3461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(297), ack => WPIPE_maxpool_output_pipe_1795_inst_req_1); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_update_completed_
      -- CP-element group 298: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1795_Update/ack
      -- 
    ack_3462_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1795_inst_ack_1, ack => convolution3D_CP_1115_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	269 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_sample_start_
      -- CP-element group 299: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Sample/$entry
      -- CP-element group 299: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Sample/req
      -- 
    req_3470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(299), ack => WPIPE_maxpool_output_pipe_1798_inst_req_0); -- 
    convolution3D_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(269) & convolution3D_CP_1115_elements(298);
      gj_convolution3D_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  transition  input  output  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (6) 
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_sample_completed_
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_update_start_
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Update/req
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Update/$entry
      -- CP-element group 300: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Sample/ack
      -- 
    ack_3471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1798_inst_ack_0, ack => convolution3D_CP_1115_elements(300)); -- 
    req_3475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(300), ack => WPIPE_maxpool_output_pipe_1798_inst_req_1); -- 
    -- CP-element group 301:  transition  input  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	302 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_update_completed_
      -- CP-element group 301: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Update/ack
      -- CP-element group 301: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1798_Update/$exit
      -- 
    ack_3476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1798_inst_ack_1, ack => convolution3D_CP_1115_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	267 
    -- CP-element group 302: 	301 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_sample_start_
      -- CP-element group 302: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Sample/$entry
      -- 
    req_3484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(302), ack => WPIPE_maxpool_output_pipe_1801_inst_req_0); -- 
    convolution3D_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(267) & convolution3D_CP_1115_elements(301);
      gj_convolution3D_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  transition  input  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (6) 
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_update_start_
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Update/req
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Sample/ack
      -- CP-element group 303: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Sample/$exit
      -- 
    ack_3485_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1801_inst_ack_0, ack => convolution3D_CP_1115_elements(303)); -- 
    req_3489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(303), ack => WPIPE_maxpool_output_pipe_1801_inst_req_1); -- 
    -- CP-element group 304:  transition  place  input  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (16) 
      -- CP-element group 304: 	 $exit
      -- CP-element group 304: 	 branch_block_stmt_441/$exit
      -- CP-element group 304: 	 branch_block_stmt_441/branch_block_stmt_441__exit__
      -- CP-element group 304: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803__exit__
      -- CP-element group 304: 	 branch_block_stmt_441/return__
      -- CP-element group 304: 	 branch_block_stmt_441/merge_stmt_1806__exit__
      -- CP-element group 304: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_update_completed_
      -- CP-element group 304: 	 branch_block_stmt_441/merge_stmt_1806_PhiReqMerge
      -- CP-element group 304: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Update/ack
      -- CP-element group 304: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/WPIPE_maxpool_output_pipe_1801_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_441/call_stmt_1695_to_assign_stmt_1803/$exit
      -- CP-element group 304: 	 branch_block_stmt_441/return___PhiReq/$entry
      -- CP-element group 304: 	 branch_block_stmt_441/return___PhiReq/$exit
      -- CP-element group 304: 	 branch_block_stmt_441/merge_stmt_1806_PhiAck/$entry
      -- CP-element group 304: 	 branch_block_stmt_441/merge_stmt_1806_PhiAck/$exit
      -- CP-element group 304: 	 branch_block_stmt_441/merge_stmt_1806_PhiAck/dummy
      -- 
    ack_3490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1801_inst_ack_1, ack => convolution3D_CP_1115_elements(304)); -- 
    -- CP-element group 305:  transition  output  delay-element  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	86 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	309 
    -- CP-element group 305:  members (5) 
      -- CP-element group 305: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_req
      -- CP-element group 305: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_757_konst_delay_trans
      -- CP-element group 305: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/$exit
      -- CP-element group 305: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/phi_stmt_751/$exit
      -- CP-element group 305: 	 branch_block_stmt_441/bbx_xnph385_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_751_req_3513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_751_req_3513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(305), ack => phi_stmt_751_req_1); -- 
    -- Element group convolution3D_CP_1115_elements(305) is a control-delay.
    cp_element_305_delay: control_delay_element  generic map(name => " 305_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(86), ack => convolution3D_CP_1115_elements(305), clk => clk, reset =>reset);
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	128 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/ra
      -- CP-element group 306: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Sample/$exit
      -- 
    ra_3533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_754_inst_ack_0, ack => convolution3D_CP_1115_elements(306)); -- 
    -- CP-element group 307:  transition  input  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	128 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/$exit
      -- CP-element group 307: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/Update/ca
      -- 
    ca_3538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_754_inst_ack_1, ack => convolution3D_CP_1115_elements(307)); -- 
    -- CP-element group 308:  join  transition  output  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (6) 
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_req
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/SplitProtocol/$exit
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/type_cast_754/$exit
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/phi_stmt_751_sources/$exit
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/phi_stmt_751/$exit
      -- CP-element group 308: 	 branch_block_stmt_441/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_751_req_3539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_751_req_3539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(308), ack => phi_stmt_751_req_0); -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(306) & convolution3D_CP_1115_elements(307);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  merge  transition  place  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	305 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	310 
    -- CP-element group 309:  members (2) 
      -- CP-element group 309: 	 branch_block_stmt_441/merge_stmt_750_PhiAck/$entry
      -- CP-element group 309: 	 branch_block_stmt_441/merge_stmt_750_PhiReqMerge
      -- 
    convolution3D_CP_1115_elements(309) <= OrReduce(convolution3D_CP_1115_elements(305) & convolution3D_CP_1115_elements(308));
    -- CP-element group 310:  fork  transition  place  input  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	309 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	87 
    -- CP-element group 310: 	88 
    -- CP-element group 310: 	90 
    -- CP-element group 310: 	91 
    -- CP-element group 310: 	94 
    -- CP-element group 310: 	98 
    -- CP-element group 310: 	102 
    -- CP-element group 310: 	106 
    -- CP-element group 310: 	110 
    -- CP-element group 310: 	114 
    -- CP-element group 310: 	118 
    -- CP-element group 310: 	122 
    -- CP-element group 310: 	125 
    -- CP-element group 310:  members (56) 
      -- CP-element group 310: 	 branch_block_stmt_441/merge_stmt_750__exit__
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913__entry__
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_resized_1
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_scaled_1
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_computed_1
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_resize_1/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_resize_1/$exit
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_resize_1/index_resize_req
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_resize_1/index_resize_ack
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_scale_1/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_scale_1/$exit
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_scale_1/scale_rename_req
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_index_scale_1/scale_rename_ack
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_update_start
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/array_obj_ref_763_final_index_sum_regn_Update/req
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_complete/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/addr_of_764_complete/req
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/RPIPE_maxpool_input_pipe_767_Sample/rr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_771_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_784_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_802_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_820_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_838_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_856_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_874_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/type_cast_892_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_update_start_
      -- CP-element group 310: 	 branch_block_stmt_441/merge_stmt_750_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/word_0/$entry
      -- CP-element group 310: 	 branch_block_stmt_441/assign_stmt_765_to_assign_stmt_913/ptr_deref_900_Update/word_access_complete/word_0/cr
      -- CP-element group 310: 	 branch_block_stmt_441/merge_stmt_750_PhiAck/phi_stmt_751_ack
      -- 
    phi_stmt_751_ack_3544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 310_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_751_ack_0, ack => convolution3D_CP_1115_elements(310)); -- 
    req_1819_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1819_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => array_obj_ref_763_index_offset_req_0); -- 
    req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => array_obj_ref_763_index_offset_req_1); -- 
    req_1839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => addr_of_764_final_reg_req_1); -- 
    rr_1848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => RPIPE_maxpool_input_pipe_767_inst_req_0); -- 
    cr_1867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_771_inst_req_1); -- 
    cr_1895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_784_inst_req_1); -- 
    cr_1923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_802_inst_req_1); -- 
    cr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_820_inst_req_1); -- 
    cr_1979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_838_inst_req_1); -- 
    cr_2007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_856_inst_req_1); -- 
    cr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_874_inst_req_1); -- 
    cr_2063_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2063_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => type_cast_892_inst_req_1); -- 
    cr_2113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(310), ack => ptr_deref_900_store_0_req_1); -- 
    -- CP-element group 311:  transition  output  delay-element  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	76 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	315 
    -- CP-element group 311:  members (5) 
      -- CP-element group 311: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_req
      -- CP-element group 311: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_951_konst_delay_trans
      -- CP-element group 311: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/$exit
      -- CP-element group 311: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/phi_stmt_945/$exit
      -- CP-element group 311: 	 branch_block_stmt_441/entry_forx_xend_PhiReq/$exit
      -- 
    phi_stmt_945_req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(311), ack => phi_stmt_945_req_1); -- 
    -- Element group convolution3D_CP_1115_elements(311) is a control-delay.
    cp_element_311_delay: control_delay_element  generic map(name => " 311_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(76), ack => convolution3D_CP_1115_elements(311), clk => clk, reset =>reset);
    -- CP-element group 312:  transition  input  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	127 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Sample/ra
      -- 
    ra_3587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_948_inst_ack_0, ack => convolution3D_CP_1115_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	127 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	314 
    -- CP-element group 313:  members (2) 
      -- CP-element group 313: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/Update/ca
      -- 
    ca_3592_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_948_inst_ack_1, ack => convolution3D_CP_1115_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: 	313 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (6) 
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/$exit
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/$exit
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_sources/type_cast_948/SplitProtocol/$exit
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/$exit
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/$exit
      -- CP-element group 314: 	 branch_block_stmt_441/forx_xcondx_xforx_xend_crit_edge_forx_xend_PhiReq/phi_stmt_945/phi_stmt_945_req
      -- 
    phi_stmt_945_req_3593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_945_req_3593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(314), ack => phi_stmt_945_req_0); -- 
    convolution3D_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(312) & convolution3D_CP_1115_elements(313);
      gj_convolution3D_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  merge  transition  place  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	311 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	316 
    -- CP-element group 315:  members (2) 
      -- CP-element group 315: 	 branch_block_stmt_441/merge_stmt_944_PhiReqMerge
      -- CP-element group 315: 	 branch_block_stmt_441/merge_stmt_944_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(315) <= OrReduce(convolution3D_CP_1115_elements(311) & convolution3D_CP_1115_elements(314));
    -- CP-element group 316:  branch  transition  place  input  output  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	315 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	129 
    -- CP-element group 316: 	130 
    -- CP-element group 316:  members (15) 
      -- CP-element group 316: 	 branch_block_stmt_441/merge_stmt_944__exit__
      -- CP-element group 316: 	 branch_block_stmt_441/assign_stmt_958_to_assign_stmt_964__entry__
      -- CP-element group 316: 	 branch_block_stmt_441/assign_stmt_958_to_assign_stmt_964__exit__
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965__entry__
      -- CP-element group 316: 	 branch_block_stmt_441/assign_stmt_958_to_assign_stmt_964/$entry
      -- CP-element group 316: 	 branch_block_stmt_441/assign_stmt_958_to_assign_stmt_964/$exit
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_dead_link/$entry
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_eval_test/$entry
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_eval_test/$exit
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_eval_test/branch_req
      -- CP-element group 316: 	 branch_block_stmt_441/R_tobool_966_place
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_if_link/$entry
      -- CP-element group 316: 	 branch_block_stmt_441/if_stmt_965_else_link/$entry
      -- CP-element group 316: 	 branch_block_stmt_441/merge_stmt_944_PhiAck/phi_stmt_945_ack
      -- CP-element group 316: 	 branch_block_stmt_441/merge_stmt_944_PhiAck/$exit
      -- 
    phi_stmt_945_ack_3598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_945_ack_0, ack => convolution3D_CP_1115_elements(316)); -- 
    branch_req_2147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(316), ack => if_stmt_965_branch_req_0); -- 
    -- CP-element group 317:  transition  output  delay-element  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	130 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (4) 
      -- CP-element group 317: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/$exit
      -- CP-element group 317: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_990_konst_delay_trans
      -- CP-element group 317: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/$exit
      -- CP-element group 317: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_req
      -- 
    phi_stmt_986_req_3621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_986_req_3621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(317), ack => phi_stmt_986_req_0); -- 
    -- Element group convolution3D_CP_1115_elements(317) is a control-delay.
    cp_element_317_delay: control_delay_element  generic map(name => " 317_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(130), ack => convolution3D_CP_1115_elements(317), clk => clk, reset =>reset);
    -- CP-element group 318:  transition  output  delay-element  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	130 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (4) 
      -- CP-element group 318: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_req
      -- CP-element group 318: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_997_konst_delay_trans
      -- CP-element group 318: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/$exit
      -- CP-element group 318: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/$exit
      -- 
    phi_stmt_993_req_3629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_993_req_3629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(318), ack => phi_stmt_993_req_0); -- 
    -- Element group convolution3D_CP_1115_elements(318) is a control-delay.
    cp_element_318_delay: control_delay_element  generic map(name => " 318_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(130), ack => convolution3D_CP_1115_elements(318), clk => clk, reset =>reset);
    -- CP-element group 319:  join  transition  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	327 
    -- CP-element group 319:  members (1) 
      -- CP-element group 319: 	 branch_block_stmt_441/bbx_xnphx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(317) & convolution3D_CP_1115_elements(318);
      gj_convolution3D_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  transition  input  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	138 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	322 
    -- CP-element group 320:  members (2) 
      -- CP-element group 320: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Sample/ra
      -- 
    ra_3649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_992_inst_ack_0, ack => convolution3D_CP_1115_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	138 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	322 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Update/$exit
      -- CP-element group 321: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/Update/ca
      -- 
    ca_3654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_992_inst_ack_1, ack => convolution3D_CP_1115_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	320 
    -- CP-element group 322: 	321 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	326 
    -- CP-element group 322:  members (5) 
      -- CP-element group 322: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/SplitProtocol/$exit
      -- CP-element group 322: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_req
      -- CP-element group 322: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/type_cast_992/$exit
      -- CP-element group 322: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/phi_stmt_986_sources/$exit
      -- CP-element group 322: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_986/$exit
      -- 
    phi_stmt_986_req_3655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_986_req_3655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(322), ack => phi_stmt_986_req_1); -- 
    convolution3D_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(320) & convolution3D_CP_1115_elements(321);
      gj_convolution3D_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	138 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Sample/ra
      -- CP-element group 323: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Sample/$exit
      -- 
    ra_3672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_0, ack => convolution3D_CP_1115_elements(323)); -- 
    -- CP-element group 324:  transition  input  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	138 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (2) 
      -- CP-element group 324: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Update/ca
      -- CP-element group 324: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/Update/$exit
      -- 
    ca_3677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_999_inst_ack_1, ack => convolution3D_CP_1115_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (5) 
      -- CP-element group 325: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/$exit
      -- CP-element group 325: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_req
      -- CP-element group 325: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/SplitProtocol/$exit
      -- CP-element group 325: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/type_cast_999/$exit
      -- CP-element group 325: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_993/phi_stmt_993_sources/$exit
      -- 
    phi_stmt_993_req_3678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_993_req_3678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(325), ack => phi_stmt_993_req_1); -- 
    convolution3D_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(323) & convolution3D_CP_1115_elements(324);
      gj_convolution3D_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	322 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	327 
    -- CP-element group 326:  members (1) 
      -- CP-element group 326: 	 branch_block_stmt_441/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(322) & convolution3D_CP_1115_elements(325);
      gj_convolution3D_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  merge  fork  transition  place  bypass 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	319 
    -- CP-element group 327: 	326 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	328 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (2) 
      -- CP-element group 327: 	 branch_block_stmt_441/merge_stmt_985_PhiReqMerge
      -- CP-element group 327: 	 branch_block_stmt_441/merge_stmt_985_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(327) <= OrReduce(convolution3D_CP_1115_elements(319) & convolution3D_CP_1115_elements(326));
    -- CP-element group 328:  transition  input  bypass 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	327 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (1) 
      -- CP-element group 328: 	 branch_block_stmt_441/merge_stmt_985_PhiAck/phi_stmt_986_ack
      -- 
    phi_stmt_986_ack_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_986_ack_0, ack => convolution3D_CP_1115_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	330 
    -- CP-element group 329:  members (1) 
      -- CP-element group 329: 	 branch_block_stmt_441/merge_stmt_985_PhiAck/phi_stmt_993_ack
      -- 
    phi_stmt_993_ack_3684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_993_ack_0, ack => convolution3D_CP_1115_elements(329)); -- 
    -- CP-element group 330:  join  fork  transition  place  output  bypass 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: 	329 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	131 
    -- CP-element group 330: 	134 
    -- CP-element group 330: 	135 
    -- CP-element group 330: 	136 
    -- CP-element group 330:  members (16) 
      -- CP-element group 330: 	 branch_block_stmt_441/merge_stmt_985__exit__
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039__entry__
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/$entry
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/RPIPE_maxpool_input_pipe_1014_Sample/rr
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_update_start_
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1018_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_update_start_
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Sample/$entry
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Sample/rr
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_441/assign_stmt_1006_to_assign_stmt_1039/type_cast_1033_Update/cr
      -- CP-element group 330: 	 branch_block_stmt_441/merge_stmt_985_PhiAck/$exit
      -- 
    rr_2172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(330), ack => RPIPE_maxpool_input_pipe_1014_inst_req_0); -- 
    cr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(330), ack => type_cast_1018_inst_req_1); -- 
    rr_2200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(330), ack => type_cast_1033_inst_req_0); -- 
    cr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(330), ack => type_cast_1033_inst_req_1); -- 
    convolution3D_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(328) & convolution3D_CP_1115_elements(329);
      gj_convolution3D_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  transition  input  bypass 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	139 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (2) 
      -- CP-element group 331: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Sample/ra
      -- 
    ra_3708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_0, ack => convolution3D_CP_1115_elements(331)); -- 
    -- CP-element group 332:  transition  input  bypass 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	139 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	333 
    -- CP-element group 332:  members (2) 
      -- CP-element group 332: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/Update/ca
      -- 
    ca_3713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_1, ack => convolution3D_CP_1115_elements(332)); -- 
    -- CP-element group 333:  join  transition  place  output  bypass 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: 	332 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	334 
    -- CP-element group 333:  members (8) 
      -- CP-element group 333: 	 branch_block_stmt_441/merge_stmt_1046_PhiReqMerge
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/SplitProtocol/$exit
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/type_cast_1050/$exit
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_sources/$exit
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/$exit
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- CP-element group 333: 	 branch_block_stmt_441/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1047/phi_stmt_1047_req
      -- CP-element group 333: 	 branch_block_stmt_441/merge_stmt_1046_PhiAck/$entry
      -- 
    phi_stmt_1047_req_3714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1047_req_3714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(333), ack => phi_stmt_1047_req_0); -- 
    convolution3D_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(331) & convolution3D_CP_1115_elements(332);
      gj_convolution3D_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	333 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	140 
    -- CP-element group 334: 	141 
    -- CP-element group 334: 	143 
    -- CP-element group 334: 	145 
    -- CP-element group 334:  members (29) 
      -- CP-element group 334: 	 branch_block_stmt_441/merge_stmt_1046__exit__
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085__entry__
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_update_start_
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_resized_1
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_scaled_1
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_computed_1
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_resize_1/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_resize_1/$exit
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_resize_1/index_resize_req
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_resize_1/index_resize_ack
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_scale_1/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_scale_1/$exit
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_scale_1/scale_rename_req
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_index_scale_1/scale_rename_ack
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_update_start
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Sample/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Sample/req
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/array_obj_ref_1079_final_index_sum_regn_Update/req
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_complete/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/addr_of_1080_complete/req
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_update_start_
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/word_0/$entry
      -- CP-element group 334: 	 branch_block_stmt_441/assign_stmt_1057_to_assign_stmt_1085/ptr_deref_1083_Update/word_access_complete/word_0/cr
      -- CP-element group 334: 	 branch_block_stmt_441/merge_stmt_1046_PhiAck/$exit
      -- CP-element group 334: 	 branch_block_stmt_441/merge_stmt_1046_PhiAck/phi_stmt_1047_ack
      -- 
    phi_stmt_1047_ack_3719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1047_ack_0, ack => convolution3D_CP_1115_elements(334)); -- 
    req_2253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(334), ack => array_obj_ref_1079_index_offset_req_0); -- 
    req_2258_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2258_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(334), ack => array_obj_ref_1079_index_offset_req_1); -- 
    req_2273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(334), ack => addr_of_1080_final_reg_req_1); -- 
    cr_2323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(334), ack => ptr_deref_1083_store_0_req_1); -- 
    -- CP-element group 335:  merge  fork  transition  place  output  bypass 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	129 
    -- CP-element group 335: 	146 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	147 
    -- CP-element group 335: 	148 
    -- CP-element group 335: 	149 
    -- CP-element group 335: 	150 
    -- CP-element group 335: 	151 
    -- CP-element group 335: 	152 
    -- CP-element group 335: 	153 
    -- CP-element group 335: 	154 
    -- CP-element group 335:  members (31) 
      -- CP-element group 335: 	 branch_block_stmt_441/merge_stmt_1087_PhiReqMerge
      -- CP-element group 335: 	 branch_block_stmt_441/merge_stmt_1087__exit__
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139__entry__
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_update_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1090_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_update_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1094_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_update_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1098_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_sample_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_update_start_
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Sample/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Sample/rr
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Update/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/assign_stmt_1091_to_assign_stmt_1139/type_cast_1102_Update/cr
      -- CP-element group 335: 	 branch_block_stmt_441/merge_stmt_1087_PhiAck/$entry
      -- CP-element group 335: 	 branch_block_stmt_441/merge_stmt_1087_PhiAck/$exit
      -- CP-element group 335: 	 branch_block_stmt_441/merge_stmt_1087_PhiAck/dummy
      -- 
    rr_2335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1090_inst_req_0); -- 
    cr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1090_inst_req_1); -- 
    rr_2349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1094_inst_req_0); -- 
    cr_2354_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2354_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1094_inst_req_1); -- 
    rr_2363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1098_inst_req_0); -- 
    cr_2368_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2368_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1098_inst_req_1); -- 
    rr_2377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1102_inst_req_0); -- 
    cr_2382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(335), ack => type_cast_1102_inst_req_1); -- 
    convolution3D_CP_1115_elements(335) <= OrReduce(convolution3D_CP_1115_elements(129) & convolution3D_CP_1115_elements(146));
    -- CP-element group 336:  transition  output  delay-element  bypass 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	170 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	340 
    -- CP-element group 336:  members (5) 
      -- CP-element group 336: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/$exit
      -- CP-element group 336: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/$exit
      -- CP-element group 336: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/$exit
      -- CP-element group 336: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1224_konst_delay_trans
      -- CP-element group 336: 	 branch_block_stmt_441/bbx_xnph_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_req
      -- 
    phi_stmt_1220_req_3753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1220_req_3753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(336), ack => phi_stmt_1220_req_0); -- 
    -- Element group convolution3D_CP_1115_elements(336) is a control-delay.
    cp_element_336_delay: control_delay_element  generic map(name => " 336_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(170), ack => convolution3D_CP_1115_elements(336), clk => clk, reset =>reset);
    -- CP-element group 337:  transition  input  bypass 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	212 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (2) 
      -- CP-element group 337: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Sample/$exit
      -- CP-element group 337: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Sample/ra
      -- 
    ra_3773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_0, ack => convolution3D_CP_1115_elements(337)); -- 
    -- CP-element group 338:  transition  input  bypass 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	212 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	339 
    -- CP-element group 338:  members (2) 
      -- CP-element group 338: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Update/$exit
      -- CP-element group 338: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/Update/ca
      -- 
    ca_3778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 338_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1226_inst_ack_1, ack => convolution3D_CP_1115_elements(338)); -- 
    -- CP-element group 339:  join  transition  output  bypass 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: 	338 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	340 
    -- CP-element group 339:  members (6) 
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/$exit
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/$exit
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/$exit
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/$exit
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_sources/type_cast_1226/SplitProtocol/$exit
      -- CP-element group 339: 	 branch_block_stmt_441/forx_xbody163_forx_xbody163_PhiReq/phi_stmt_1220/phi_stmt_1220_req
      -- 
    phi_stmt_1220_req_3779_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1220_req_3779_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(339), ack => phi_stmt_1220_req_1); -- 
    convolution3D_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(337) & convolution3D_CP_1115_elements(338);
      gj_convolution3D_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  merge  transition  place  bypass 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	336 
    -- CP-element group 340: 	339 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	341 
    -- CP-element group 340:  members (2) 
      -- CP-element group 340: 	 branch_block_stmt_441/merge_stmt_1219_PhiReqMerge
      -- CP-element group 340: 	 branch_block_stmt_441/merge_stmt_1219_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(340) <= OrReduce(convolution3D_CP_1115_elements(336) & convolution3D_CP_1115_elements(339));
    -- CP-element group 341:  fork  transition  place  input  output  bypass 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	340 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	171 
    -- CP-element group 341: 	172 
    -- CP-element group 341: 	174 
    -- CP-element group 341: 	175 
    -- CP-element group 341: 	178 
    -- CP-element group 341: 	182 
    -- CP-element group 341: 	186 
    -- CP-element group 341: 	190 
    -- CP-element group 341: 	194 
    -- CP-element group 341: 	198 
    -- CP-element group 341: 	202 
    -- CP-element group 341: 	206 
    -- CP-element group 341: 	209 
    -- CP-element group 341:  members (56) 
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_resize_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_scale_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_scaled_1
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_scale_1/scale_rename_ack
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_scale_1/scale_rename_req
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_resized_1
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_scale_1/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_computed_1
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_resize_1/$exit
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_resize_1/index_resize_req
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/RPIPE_maxpool_input_pipe_1236_Sample/rr
      -- CP-element group 341: 	 branch_block_stmt_441/merge_stmt_1219__exit__
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382__entry__
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_update_start
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Sample/req
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_complete/req
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1253_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_index_resize_1/index_resize_ack
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/addr_of_1233_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1343_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1325_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1289_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1307_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Update/req
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1240_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1271_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/array_obj_ref_1232_final_index_sum_regn_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/type_cast_1361_Update/cr
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_update_start_
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/word_0/$entry
      -- CP-element group 341: 	 branch_block_stmt_441/assign_stmt_1234_to_assign_stmt_1382/ptr_deref_1369_Update/word_access_complete/word_0/cr
      -- CP-element group 341: 	 branch_block_stmt_441/merge_stmt_1219_PhiAck/$exit
      -- CP-element group 341: 	 branch_block_stmt_441/merge_stmt_1219_PhiAck/phi_stmt_1220_ack
      -- 
    phi_stmt_1220_ack_3784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1220_ack_0, ack => convolution3D_CP_1115_elements(341)); -- 
    cr_2593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1253_inst_req_1); -- 
    rr_2546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => RPIPE_maxpool_input_pipe_1236_inst_req_0); -- 
    req_2517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => array_obj_ref_1232_index_offset_req_0); -- 
    cr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1325_inst_req_1); -- 
    req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => addr_of_1233_final_reg_req_1); -- 
    cr_2677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1307_inst_req_1); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1343_inst_req_1); -- 
    cr_2621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1271_inst_req_1); -- 
    cr_2565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1240_inst_req_1); -- 
    cr_2649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1289_inst_req_1); -- 
    req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => array_obj_ref_1232_index_offset_req_1); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => type_cast_1361_inst_req_1); -- 
    cr_2811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(341), ack => ptr_deref_1369_store_0_req_1); -- 
    -- CP-element group 342:  transition  input  bypass 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	211 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (2) 
      -- CP-element group 342: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Sample/$exit
      -- CP-element group 342: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Sample/ra
      -- 
    ra_3816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 342_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_0, ack => convolution3D_CP_1115_elements(342)); -- 
    -- CP-element group 343:  transition  input  bypass 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	211 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	344 
    -- CP-element group 343:  members (2) 
      -- CP-element group 343: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Update/$exit
      -- CP-element group 343: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/Update/ca
      -- 
    ca_3821_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1417_inst_ack_1, ack => convolution3D_CP_1115_elements(343)); -- 
    -- CP-element group 344:  join  transition  output  bypass 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	343 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	346 
    -- CP-element group 344:  members (6) 
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/$exit
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/$exit
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/$exit
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/$exit
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1417/SplitProtocol/$exit
      -- CP-element group 344: 	 branch_block_stmt_441/forx_xcond156x_xforx_xend215_crit_edge_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_req
      -- 
    phi_stmt_1414_req_3822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1414_req_3822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(344), ack => phi_stmt_1414_req_0); -- 
    convolution3D_cp_element_group_344: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_344"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(342) & convolution3D_CP_1115_elements(343);
      gj_convolution3D_cp_element_group_344 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(344), clk => clk, reset => reset); --
    end block;
    -- CP-element group 345:  transition  output  delay-element  bypass 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	157 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (5) 
      -- CP-element group 345: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/$exit
      -- CP-element group 345: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/$exit
      -- CP-element group 345: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/$exit
      -- CP-element group 345: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_sources/type_cast_1420_konst_delay_trans
      -- CP-element group 345: 	 branch_block_stmt_441/ifx_xend_forx_xend215_PhiReq/phi_stmt_1414/phi_stmt_1414_req
      -- 
    phi_stmt_1414_req_3833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1414_req_3833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(345), ack => phi_stmt_1414_req_1); -- 
    -- Element group convolution3D_CP_1115_elements(345) is a control-delay.
    cp_element_345_delay: control_delay_element  generic map(name => " 345_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(157), ack => convolution3D_CP_1115_elements(345), clk => clk, reset =>reset);
    -- CP-element group 346:  merge  transition  place  bypass 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	344 
    -- CP-element group 346: 	345 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (2) 
      -- CP-element group 346: 	 branch_block_stmt_441/merge_stmt_1413_PhiReqMerge
      -- CP-element group 346: 	 branch_block_stmt_441/merge_stmt_1413_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(346) <= OrReduce(convolution3D_CP_1115_elements(344) & convolution3D_CP_1115_elements(345));
    -- CP-element group 347:  branch  transition  place  input  output  bypass 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	213 
    -- CP-element group 347: 	214 
    -- CP-element group 347:  members (15) 
      -- CP-element group 347: 	 branch_block_stmt_441/R_tobool218_1435_place
      -- CP-element group 347: 	 branch_block_stmt_441/merge_stmt_1413__exit__
      -- CP-element group 347: 	 branch_block_stmt_441/assign_stmt_1427_to_assign_stmt_1433__entry__
      -- CP-element group 347: 	 branch_block_stmt_441/assign_stmt_1427_to_assign_stmt_1433__exit__
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434__entry__
      -- CP-element group 347: 	 branch_block_stmt_441/assign_stmt_1427_to_assign_stmt_1433/$entry
      -- CP-element group 347: 	 branch_block_stmt_441/assign_stmt_1427_to_assign_stmt_1433/$exit
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_dead_link/$entry
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_eval_test/$entry
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_eval_test/$exit
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_eval_test/branch_req
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_if_link/$entry
      -- CP-element group 347: 	 branch_block_stmt_441/if_stmt_1434_else_link/$entry
      -- CP-element group 347: 	 branch_block_stmt_441/merge_stmt_1413_PhiAck/$exit
      -- CP-element group 347: 	 branch_block_stmt_441/merge_stmt_1413_PhiAck/phi_stmt_1414_ack
      -- 
    phi_stmt_1414_ack_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1414_ack_0, ack => convolution3D_CP_1115_elements(347)); -- 
    branch_req_2845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(347), ack => if_stmt_1434_branch_req_0); -- 
    -- CP-element group 348:  transition  output  delay-element  bypass 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	216 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	350 
    -- CP-element group 348:  members (4) 
      -- CP-element group 348: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/$exit
      -- CP-element group 348: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/$exit
      -- CP-element group 348: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1463_konst_delay_trans
      -- CP-element group 348: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_req
      -- 
    phi_stmt_1459_req_3861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1459_req_3861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(348), ack => phi_stmt_1459_req_0); -- 
    -- Element group convolution3D_CP_1115_elements(348) is a control-delay.
    cp_element_348_delay: control_delay_element  generic map(name => " 348_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(216), ack => convolution3D_CP_1115_elements(348), clk => clk, reset =>reset);
    -- CP-element group 349:  transition  output  delay-element  bypass 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	216 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	350 
    -- CP-element group 349:  members (4) 
      -- CP-element group 349: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/$exit
      -- CP-element group 349: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$exit
      -- CP-element group 349: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1470_konst_delay_trans
      -- CP-element group 349: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_req
      -- 
    phi_stmt_1466_req_3869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1466_req_3869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(349), ack => phi_stmt_1466_req_0); -- 
    -- Element group convolution3D_CP_1115_elements(349) is a control-delay.
    cp_element_349_delay: control_delay_element  generic map(name => " 349_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(216), ack => convolution3D_CP_1115_elements(349), clk => clk, reset =>reset);
    -- CP-element group 350:  join  transition  bypass 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	348 
    -- CP-element group 350: 	349 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	358 
    -- CP-element group 350:  members (1) 
      -- CP-element group 350: 	 branch_block_stmt_441/bbx_xnphx_xi356_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(348) & convolution3D_CP_1115_elements(349);
      gj_convolution3D_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  transition  input  bypass 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	224 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (2) 
      -- CP-element group 351: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Sample/ra
      -- 
    ra_3889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1465_inst_ack_0, ack => convolution3D_CP_1115_elements(351)); -- 
    -- CP-element group 352:  transition  input  bypass 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	224 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	353 
    -- CP-element group 352:  members (2) 
      -- CP-element group 352: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/Update/ca
      -- 
    ca_3894_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1465_inst_ack_1, ack => convolution3D_CP_1115_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: 	352 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	357 
    -- CP-element group 353:  members (5) 
      -- CP-element group 353: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/$exit
      -- CP-element group 353: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/$exit
      -- CP-element group 353: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/$exit
      -- CP-element group 353: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_sources/type_cast_1465/SplitProtocol/$exit
      -- CP-element group 353: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1459/phi_stmt_1459_req
      -- 
    phi_stmt_1459_req_3895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1459_req_3895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(353), ack => phi_stmt_1459_req_1); -- 
    convolution3D_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(351) & convolution3D_CP_1115_elements(352);
      gj_convolution3D_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  transition  input  bypass 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	224 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (2) 
      -- CP-element group 354: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Sample/$exit
      -- CP-element group 354: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Sample/ra
      -- 
    ra_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_0, ack => convolution3D_CP_1115_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	224 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (2) 
      -- CP-element group 355: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Update/$exit
      -- CP-element group 355: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/Update/ca
      -- 
    ca_3917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1472_inst_ack_1, ack => convolution3D_CP_1115_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: 	355 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	357 
    -- CP-element group 356:  members (5) 
      -- CP-element group 356: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/$exit
      -- CP-element group 356: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$exit
      -- CP-element group 356: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/$exit
      -- CP-element group 356: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472/SplitProtocol/$exit
      -- CP-element group 356: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/phi_stmt_1466/phi_stmt_1466_req
      -- 
    phi_stmt_1466_req_3918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1466_req_3918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(356), ack => phi_stmt_1466_req_1); -- 
    convolution3D_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(354) & convolution3D_CP_1115_elements(355);
      gj_convolution3D_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  join  transition  bypass 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	353 
    -- CP-element group 357: 	356 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	358 
    -- CP-element group 357:  members (1) 
      -- CP-element group 357: 	 branch_block_stmt_441/forx_xbodyx_xi365_forx_xbodyx_xi365_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(353) & convolution3D_CP_1115_elements(356);
      gj_convolution3D_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  merge  fork  transition  place  bypass 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	350 
    -- CP-element group 358: 	357 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	359 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (2) 
      -- CP-element group 358: 	 branch_block_stmt_441/merge_stmt_1458_PhiReqMerge
      -- CP-element group 358: 	 branch_block_stmt_441/merge_stmt_1458_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(358) <= OrReduce(convolution3D_CP_1115_elements(350) & convolution3D_CP_1115_elements(357));
    -- CP-element group 359:  transition  input  bypass 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	358 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (1) 
      -- CP-element group 359: 	 branch_block_stmt_441/merge_stmt_1458_PhiAck/phi_stmt_1459_ack
      -- 
    phi_stmt_1459_ack_3923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1459_ack_0, ack => convolution3D_CP_1115_elements(359)); -- 
    -- CP-element group 360:  transition  input  bypass 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	361 
    -- CP-element group 360:  members (1) 
      -- CP-element group 360: 	 branch_block_stmt_441/merge_stmt_1458_PhiAck/phi_stmt_1466_ack
      -- 
    phi_stmt_1466_ack_3924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1466_ack_0, ack => convolution3D_CP_1115_elements(360)); -- 
    -- CP-element group 361:  join  fork  transition  place  output  bypass 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: 	360 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	217 
    -- CP-element group 361: 	220 
    -- CP-element group 361: 	221 
    -- CP-element group 361: 	222 
    -- CP-element group 361:  members (16) 
      -- CP-element group 361: 	 branch_block_stmt_441/merge_stmt_1458__exit__
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512__entry__
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/$entry
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/RPIPE_maxpool_input_pipe_1487_Sample/rr
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_update_start_
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1491_Update/cr
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_update_start_
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Sample/rr
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Update/$entry
      -- CP-element group 361: 	 branch_block_stmt_441/assign_stmt_1479_to_assign_stmt_1512/type_cast_1506_Update/cr
      -- CP-element group 361: 	 branch_block_stmt_441/merge_stmt_1458_PhiAck/$exit
      -- 
    rr_2884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(361), ack => RPIPE_maxpool_input_pipe_1487_inst_req_0); -- 
    cr_2903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(361), ack => type_cast_1491_inst_req_1); -- 
    rr_2912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(361), ack => type_cast_1506_inst_req_0); -- 
    cr_2917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(361), ack => type_cast_1506_inst_req_1); -- 
    convolution3D_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(359) & convolution3D_CP_1115_elements(360);
      gj_convolution3D_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  transition  input  bypass 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	225 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (2) 
      -- CP-element group 362: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Sample/$exit
      -- CP-element group 362: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Sample/ra
      -- 
    ra_3948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_0, ack => convolution3D_CP_1115_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	225 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (2) 
      -- CP-element group 363: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/Update/ca
      -- 
    ca_3953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1523_inst_ack_1, ack => convolution3D_CP_1115_elements(363)); -- 
    -- CP-element group 364:  join  transition  place  output  bypass 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: 	363 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (8) 
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/$exit
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/$exit
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/$exit
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/$exit
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_sources/type_cast_1523/SplitProtocol/$exit
      -- CP-element group 364: 	 branch_block_stmt_441/forx_xbodyx_xi365_getRemainingElementsx_xexit373_PhiReq/phi_stmt_1520/phi_stmt_1520_req
      -- CP-element group 364: 	 branch_block_stmt_441/merge_stmt_1519_PhiReqMerge
      -- CP-element group 364: 	 branch_block_stmt_441/merge_stmt_1519_PhiAck/$entry
      -- 
    phi_stmt_1520_req_3954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1520_req_3954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(364), ack => phi_stmt_1520_req_0); -- 
    convolution3D_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(362) & convolution3D_CP_1115_elements(363);
      gj_convolution3D_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	226 
    -- CP-element group 365: 	227 
    -- CP-element group 365: 	229 
    -- CP-element group 365: 	231 
    -- CP-element group 365:  members (29) 
      -- CP-element group 365: 	 branch_block_stmt_441/merge_stmt_1519__exit__
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558__entry__
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_update_start_
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_resized_1
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_scaled_1
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_computed_1
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_resize_1/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_resize_1/$exit
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_resize_1/index_resize_req
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_resize_1/index_resize_ack
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_scale_1/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_scale_1/$exit
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_scale_1/scale_rename_req
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_index_scale_1/scale_rename_ack
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_update_start
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Sample/req
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/array_obj_ref_1552_final_index_sum_regn_Update/req
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_complete/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/addr_of_1553_complete/req
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_update_start_
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/word_0/$entry
      -- CP-element group 365: 	 branch_block_stmt_441/assign_stmt_1530_to_assign_stmt_1558/ptr_deref_1556_Update/word_access_complete/word_0/cr
      -- CP-element group 365: 	 branch_block_stmt_441/merge_stmt_1519_PhiAck/$exit
      -- CP-element group 365: 	 branch_block_stmt_441/merge_stmt_1519_PhiAck/phi_stmt_1520_ack
      -- 
    phi_stmt_1520_ack_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1520_ack_0, ack => convolution3D_CP_1115_elements(365)); -- 
    req_2965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(365), ack => array_obj_ref_1552_index_offset_req_0); -- 
    req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(365), ack => array_obj_ref_1552_index_offset_req_1); -- 
    req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(365), ack => addr_of_1553_final_reg_req_1); -- 
    cr_3035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(365), ack => ptr_deref_1556_store_0_req_1); -- 
    -- CP-element group 366:  merge  fork  transition  place  output  bypass 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	213 
    -- CP-element group 366: 	232 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	233 
    -- CP-element group 366: 	234 
    -- CP-element group 366:  members (13) 
      -- CP-element group 366: 	 branch_block_stmt_441/merge_stmt_1560__exit__
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563__entry__
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/$entry
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_update_start_
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Sample/crr
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_441/call_stmt_1563/call_stmt_1563_Update/ccr
      -- CP-element group 366: 	 branch_block_stmt_441/merge_stmt_1560_PhiReqMerge
      -- CP-element group 366: 	 branch_block_stmt_441/merge_stmt_1560_PhiAck/$entry
      -- CP-element group 366: 	 branch_block_stmt_441/merge_stmt_1560_PhiAck/$exit
      -- CP-element group 366: 	 branch_block_stmt_441/merge_stmt_1560_PhiAck/dummy
      -- 
    crr_3047_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3047_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(366), ack => call_stmt_1563_call_req_0); -- 
    ccr_3052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(366), ack => call_stmt_1563_call_req_1); -- 
    convolution3D_CP_1115_elements(366) <= OrReduce(convolution3D_CP_1115_elements(213) & convolution3D_CP_1115_elements(232));
    -- CP-element group 367:  transition  output  delay-element  bypass 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	247 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	371 
    -- CP-element group 367:  members (5) 
      -- CP-element group 367: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/$exit
      -- CP-element group 367: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/$exit
      -- CP-element group 367: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/$exit
      -- CP-element group 367: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1640_konst_delay_trans
      -- CP-element group 367: 	 branch_block_stmt_441/ifx_xend227_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_req
      -- 
    phi_stmt_1634_req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1634_req_3981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(367), ack => phi_stmt_1634_req_1); -- 
    -- Element group convolution3D_CP_1115_elements(367) is a control-delay.
    cp_element_367_delay: control_delay_element  generic map(name => " 367_delay", delay_value => 1)  port map(req => convolution3D_CP_1115_elements(247), ack => convolution3D_CP_1115_elements(367), clk => clk, reset =>reset);
    -- CP-element group 368:  transition  input  bypass 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	259 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	370 
    -- CP-element group 368:  members (2) 
      -- CP-element group 368: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Sample/ra
      -- 
    ra_4001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1637_inst_ack_0, ack => convolution3D_CP_1115_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	259 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	370 
    -- CP-element group 369:  members (2) 
      -- CP-element group 369: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/Update/ca
      -- 
    ca_4006_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1637_inst_ack_1, ack => convolution3D_CP_1115_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	368 
    -- CP-element group 370: 	369 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	371 
    -- CP-element group 370:  members (6) 
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/$exit
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/$exit
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/$exit
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_sources/type_cast_1637/SplitProtocol/$exit
      -- CP-element group 370: 	 branch_block_stmt_441/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1634/phi_stmt_1634_req
      -- 
    phi_stmt_1634_req_4007_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1634_req_4007_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(370), ack => phi_stmt_1634_req_0); -- 
    convolution3D_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_1115_elements(368) & convolution3D_CP_1115_elements(369);
      gj_convolution3D_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_1115_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  merge  transition  place  bypass 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	367 
    -- CP-element group 371: 	370 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	372 
    -- CP-element group 371:  members (2) 
      -- CP-element group 371: 	 branch_block_stmt_441/merge_stmt_1633_PhiReqMerge
      -- CP-element group 371: 	 branch_block_stmt_441/merge_stmt_1633_PhiAck/$entry
      -- 
    convolution3D_CP_1115_elements(371) <= OrReduce(convolution3D_CP_1115_elements(367) & convolution3D_CP_1115_elements(370));
    -- CP-element group 372:  fork  transition  place  input  output  bypass 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	371 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	248 
    -- CP-element group 372: 	249 
    -- CP-element group 372: 	250 
    -- CP-element group 372: 	251 
    -- CP-element group 372: 	254 
    -- CP-element group 372: 	255 
    -- CP-element group 372: 	256 
    -- CP-element group 372:  members (26) 
      -- CP-element group 372: 	 branch_block_stmt_441/merge_stmt_1633__exit__
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680__entry__
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_update_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Sample/rr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1654_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_update_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Sample/rr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/type_cast_1658_Update/cr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_update_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1662_Update/ccr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_sample_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_update_start_
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Sample/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Sample/crr
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Update/$entry
      -- CP-element group 372: 	 branch_block_stmt_441/assign_stmt_1646_to_assign_stmt_1680/call_stmt_1669_Update/ccr
      -- CP-element group 372: 	 branch_block_stmt_441/merge_stmt_1633_PhiAck/$exit
      -- CP-element group 372: 	 branch_block_stmt_441/merge_stmt_1633_PhiAck/phi_stmt_1634_ack
      -- 
    phi_stmt_1634_ack_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1634_ack_0, ack => convolution3D_CP_1115_elements(372)); -- 
    rr_3151_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3151_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => type_cast_1654_inst_req_0); -- 
    cr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => type_cast_1654_inst_req_1); -- 
    rr_3165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => type_cast_1658_inst_req_0); -- 
    cr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => type_cast_1658_inst_req_1); -- 
    ccr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => call_stmt_1662_call_req_1); -- 
    crr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => call_stmt_1669_call_req_0); -- 
    ccr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_1115_elements(372), ack => call_stmt_1669_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i64_i64_1131_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_1409_wire : std_logic_vector(63 downto 0);
    signal ASHR_i64_i64_940_wire : std_logic_vector(63 downto 0);
    signal Bx_xnot_1057 : std_logic_vector(63 downto 0);
    signal R_indvar412_1231_resized : std_logic_vector(13 downto 0);
    signal R_indvar412_1231_scaled : std_logic_vector(13 downto 0);
    signal R_indvar426_762_resized : std_logic_vector(13 downto 0);
    signal R_indvar426_762_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1078_resized : std_logic_vector(13 downto 0);
    signal R_ix_x0x_xlcssa_1078_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1551_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1551_scaled : std_logic_vector(13 downto 0);
    signal add102_808 : std_logic_vector(63 downto 0);
    signal add108_826 : std_logic_vector(63 downto 0);
    signal add114_844 : std_logic_vector(63 downto 0);
    signal add120_862 : std_logic_vector(63 downto 0);
    signal add1216x_xi370_1536 : std_logic_vector(63 downto 0);
    signal add1216x_xi_1063 : std_logic_vector(63 downto 0);
    signal add126_880 : std_logic_vector(63 downto 0);
    signal add132_898 : std_logic_vector(63 downto 0);
    signal add13_492 : std_logic_vector(15 downto 0);
    signal add171_1259 : std_logic_vector(63 downto 0);
    signal add177_1277 : std_logic_vector(63 downto 0);
    signal add183_1295 : std_logic_vector(63 downto 0);
    signal add189_1313 : std_logic_vector(63 downto 0);
    signal add195_1331 : std_logic_vector(63 downto 0);
    signal add201_1349 : std_logic_vector(63 downto 0);
    signal add207_1367 : std_logic_vector(63 downto 0);
    signal add23_517 : std_logic_vector(15 downto 0);
    signal add33_542 : std_logic_vector(15 downto 0);
    signal add43_567 : std_logic_vector(15 downto 0);
    signal add53_592 : std_logic_vector(15 downto 0);
    signal add63_617 : std_logic_vector(15 downto 0);
    signal add73_642 : std_logic_vector(15 downto 0);
    signal add96_790 : std_logic_vector(63 downto 0);
    signal add_467 : std_logic_vector(31 downto 0);
    signal addx_xi361_1497 : std_logic_vector(63 downto 0);
    signal addx_xi_1024 : std_logic_vector(63 downto 0);
    signal and217_1427 : std_logic_vector(63 downto 0);
    signal and_958 : std_logic_vector(63 downto 0);
    signal array_obj_ref_1079_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1079_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1232_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1552_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_763_root_address : std_logic_vector(13 downto 0);
    signal arrayidx143_1081 : std_logic_vector(31 downto 0);
    signal arrayidx211_1234 : std_logic_vector(31 downto 0);
    signal arrayidx226_1554 : std_logic_vector(31 downto 0);
    signal arrayidx_765 : std_logic_vector(31 downto 0);
    signal call105_817 : std_logic_vector(7 downto 0);
    signal call111_835 : std_logic_vector(7 downto 0);
    signal call117_853 : std_logic_vector(7 downto 0);
    signal call11_483 : std_logic_vector(7 downto 0);
    signal call123_871 : std_logic_vector(7 downto 0);
    signal call129_889 : std_logic_vector(7 downto 0);
    signal call164_1237 : std_logic_vector(7 downto 0);
    signal call168_1250 : std_logic_vector(7 downto 0);
    signal call16_495 : std_logic_vector(7 downto 0);
    signal call174_1268 : std_logic_vector(7 downto 0);
    signal call180_1286 : std_logic_vector(7 downto 0);
    signal call186_1304 : std_logic_vector(7 downto 0);
    signal call192_1322 : std_logic_vector(7 downto 0);
    signal call198_1340 : std_logic_vector(7 downto 0);
    signal call204_1358 : std_logic_vector(7 downto 0);
    signal call21_508 : std_logic_vector(7 downto 0);
    signal call229_1563 : std_logic_vector(63 downto 0);
    signal call26_520 : std_logic_vector(7 downto 0);
    signal call284_1695 : std_logic_vector(63 downto 0);
    signal call2_458 : std_logic_vector(7 downto 0);
    signal call31_533 : std_logic_vector(7 downto 0);
    signal call36_545 : std_logic_vector(7 downto 0);
    signal call41_558 : std_logic_vector(7 downto 0);
    signal call46_570 : std_logic_vector(7 downto 0);
    signal call51_583 : std_logic_vector(7 downto 0);
    signal call56_595 : std_logic_vector(7 downto 0);
    signal call61_608 : std_logic_vector(7 downto 0);
    signal call66_620 : std_logic_vector(7 downto 0);
    signal call6_470 : std_logic_vector(7 downto 0);
    signal call71_633 : std_logic_vector(7 downto 0);
    signal call89_768 : std_logic_vector(7 downto 0);
    signal call93_781 : std_logic_vector(7 downto 0);
    signal call99_799 : std_logic_vector(7 downto 0);
    signal call_445 : std_logic_vector(7 downto 0);
    signal callx_xi359_1488 : std_logic_vector(7 downto 0);
    signal callx_xi_1015 : std_logic_vector(7 downto 0);
    signal cmp161379_1139 : std_logic_vector(0 downto 0);
    signal cmp383_672 : std_logic_vector(0 downto 0);
    signal cmpx_xi364_1512 : std_logic_vector(0 downto 0);
    signal cmpx_xi_1039 : std_logic_vector(0 downto 0);
    signal conv101_803 : std_logic_vector(63 downto 0);
    signal conv107_821 : std_logic_vector(63 downto 0);
    signal conv113_839 : std_logic_vector(63 downto 0);
    signal conv119_857 : std_logic_vector(63 downto 0);
    signal conv125_875 : std_logic_vector(63 downto 0);
    signal conv12_487 : std_logic_vector(15 downto 0);
    signal conv131_893 : std_logic_vector(63 downto 0);
    signal conv145_1091 : std_logic_vector(63 downto 0);
    signal conv147_1095 : std_logic_vector(63 downto 0);
    signal conv150_1099 : std_logic_vector(63 downto 0);
    signal conv153_1103 : std_logic_vector(63 downto 0);
    signal conv155_1133 : std_logic_vector(63 downto 0);
    signal conv165_1241 : std_logic_vector(63 downto 0);
    signal conv170_1254 : std_logic_vector(63 downto 0);
    signal conv176_1272 : std_logic_vector(63 downto 0);
    signal conv182_1290 : std_logic_vector(63 downto 0);
    signal conv188_1308 : std_logic_vector(63 downto 0);
    signal conv194_1326 : std_logic_vector(63 downto 0);
    signal conv19_499 : std_logic_vector(15 downto 0);
    signal conv1_449 : std_logic_vector(31 downto 0);
    signal conv200_1344 : std_logic_vector(63 downto 0);
    signal conv206_1362 : std_logic_vector(63 downto 0);
    signal conv22_512 : std_logic_vector(15 downto 0);
    signal conv230_1692 : std_logic_vector(63 downto 0);
    signal conv255_1655 : std_logic_vector(63 downto 0);
    signal conv261_1659 : std_logic_vector(63 downto 0);
    signal conv285_1700 : std_logic_vector(63 downto 0);
    signal conv293_1709 : std_logic_vector(7 downto 0);
    signal conv299_1719 : std_logic_vector(7 downto 0);
    signal conv29_524 : std_logic_vector(15 downto 0);
    signal conv2x_xi354_1450 : std_logic_vector(31 downto 0);
    signal conv2x_xi_977 : std_logic_vector(31 downto 0);
    signal conv305_1729 : std_logic_vector(7 downto 0);
    signal conv311_1739 : std_logic_vector(7 downto 0);
    signal conv317_1749 : std_logic_vector(7 downto 0);
    signal conv323_1759 : std_logic_vector(7 downto 0);
    signal conv329_1769 : std_logic_vector(7 downto 0);
    signal conv32_537 : std_logic_vector(15 downto 0);
    signal conv335_1779 : std_logic_vector(7 downto 0);
    signal conv39_549 : std_logic_vector(15 downto 0);
    signal conv3_462 : std_logic_vector(31 downto 0);
    signal conv42_562 : std_logic_vector(15 downto 0);
    signal conv49_574 : std_logic_vector(15 downto 0);
    signal conv52_587 : std_logic_vector(15 downto 0);
    signal conv59_599 : std_logic_vector(15 downto 0);
    signal conv5x_xi360_1492 : std_logic_vector(63 downto 0);
    signal conv5x_xi_1019 : std_logic_vector(63 downto 0);
    signal conv62_612 : std_logic_vector(15 downto 0);
    signal conv69_624 : std_logic_vector(15 downto 0);
    signal conv72_637 : std_logic_vector(15 downto 0);
    signal conv79_646 : std_logic_vector(31 downto 0);
    signal conv81_650 : std_logic_vector(31 downto 0);
    signal conv83_666 : std_logic_vector(63 downto 0);
    signal conv90_772 : std_logic_vector(63 downto 0);
    signal conv95_785 : std_logic_vector(63 downto 0);
    signal conv9_474 : std_logic_vector(15 downto 0);
    signal convx_xi363_1507 : std_logic_vector(31 downto 0);
    signal convx_xi_1034 : std_logic_vector(31 downto 0);
    signal elementx_x021x_xi358_1466 : std_logic_vector(63 downto 0);
    signal elementx_x021x_xi_993 : std_logic_vector(63 downto 0);
    signal exitcond32_913 : std_logic_vector(0 downto 0);
    signal exitcond5_1680 : std_logic_vector(0 downto 0);
    signal exitcond_1382 : std_logic_vector(0 downto 0);
    signal iNsTr_35_1012 : std_logic_vector(15 downto 0);
    signal iNsTr_57_1446 : std_logic_vector(63 downto 0);
    signal iNsTr_65_1485 : std_logic_vector(15 downto 0);
    signal iNsTr_87_1530 : std_logic_vector(63 downto 0);
    signal indvar412_1220 : std_logic_vector(63 downto 0);
    signal indvar426_751 : std_logic_vector(63 downto 0);
    signal indvar_1634 : std_logic_vector(31 downto 0);
    signal indvarx_xnext413_1377 : std_logic_vector(63 downto 0);
    signal indvarx_xnext427_908 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1675 : std_logic_vector(31 downto 0);
    signal ix_x0x_xlcssa_945 : std_logic_vector(63 downto 0);
    signal ix_x1x_xlcssa_1414 : std_logic_vector(63 downto 0);
    signal mul148_1108 : std_logic_vector(63 downto 0);
    signal mul151_1113 : std_logic_vector(63 downto 0);
    signal mul154_1118 : std_logic_vector(63 downto 0);
    signal mul236_1569 : std_logic_vector(15 downto 0);
    signal mul249_1574 : std_logic_vector(15 downto 0);
    signal mul254_1646 : std_logic_vector(31 downto 0);
    signal mul260_1651 : std_logic_vector(31 downto 0);
    signal mul82_660 : std_logic_vector(31 downto 0);
    signal mul_655 : std_logic_vector(31 downto 0);
    signal nx_x022x_xi357_1459 : std_logic_vector(15 downto 0);
    signal nx_x022x_xi_986 : std_logic_vector(15 downto 0);
    signal phitmp387_1411 : std_logic_vector(63 downto 0);
    signal phitmp_942 : std_logic_vector(63 downto 0);
    signal ptr_deref_1083_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1083_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1083_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1083_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1083_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1083_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1369_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1369_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1369_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1369_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1369_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1369_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1556_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1556_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1556_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1556_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1556_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1556_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_900_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_900_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_900_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_900_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_900_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_900_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext_1124 : std_logic_vector(63 downto 0);
    signal sh_promx_xi371_1542 : std_logic_vector(63 downto 0);
    signal sh_promx_xi_1069 : std_logic_vector(63 downto 0);
    signal shl104_814 : std_logic_vector(63 downto 0);
    signal shl10_480 : std_logic_vector(15 downto 0);
    signal shl110_832 : std_logic_vector(63 downto 0);
    signal shl116_850 : std_logic_vector(63 downto 0);
    signal shl122_868 : std_logic_vector(63 downto 0);
    signal shl128_886 : std_logic_vector(63 downto 0);
    signal shl14x_xi372_1547 : std_logic_vector(63 downto 0);
    signal shl14x_xi_1074 : std_logic_vector(63 downto 0);
    signal shl167_1247 : std_logic_vector(63 downto 0);
    signal shl173_1265 : std_logic_vector(63 downto 0);
    signal shl179_1283 : std_logic_vector(63 downto 0);
    signal shl185_1301 : std_logic_vector(63 downto 0);
    signal shl191_1319 : std_logic_vector(63 downto 0);
    signal shl197_1337 : std_logic_vector(63 downto 0);
    signal shl203_1355 : std_logic_vector(63 downto 0);
    signal shl20_505 : std_logic_vector(15 downto 0);
    signal shl30_530 : std_logic_vector(15 downto 0);
    signal shl40_555 : std_logic_vector(15 downto 0);
    signal shl50_580 : std_logic_vector(15 downto 0);
    signal shl60_605 : std_logic_vector(15 downto 0);
    signal shl70_630 : std_logic_vector(15 downto 0);
    signal shl8x_xi362_1503 : std_logic_vector(63 downto 0);
    signal shl8x_xi362x_xlcssa_1520 : std_logic_vector(63 downto 0);
    signal shl8x_xi_1030 : std_logic_vector(63 downto 0);
    signal shl8x_xix_xlcssa_1047 : std_logic_vector(63 downto 0);
    signal shl92_778 : std_logic_vector(63 downto 0);
    signal shl98_796 : std_logic_vector(63 downto 0);
    signal shl_455 : std_logic_vector(31 downto 0);
    signal shlx_xi355_1456 : std_logic_vector(31 downto 0);
    signal shlx_xi_983 : std_logic_vector(31 downto 0);
    signal shr296_1715 : std_logic_vector(63 downto 0);
    signal shr302_1725 : std_logic_vector(63 downto 0);
    signal shr308_1735 : std_logic_vector(63 downto 0);
    signal shr314_1745 : std_logic_vector(63 downto 0);
    signal shr320_1755 : std_logic_vector(63 downto 0);
    signal shr326_1765 : std_logic_vector(63 downto 0);
    signal shr332_1775 : std_logic_vector(63 downto 0);
    signal sub269_1597 : std_logic_vector(15 downto 0);
    signal sub289_1705 : std_logic_vector(63 downto 0);
    signal sub_1591 : std_logic_vector(15 downto 0);
    signal tmp12_1162 : std_logic_vector(63 downto 0);
    signal tmp13_1166 : std_logic_vector(63 downto 0);
    signal tmp14_1171 : std_logic_vector(63 downto 0);
    signal tmp15_1175 : std_logic_vector(63 downto 0);
    signal tmp16_1180 : std_logic_vector(63 downto 0);
    signal tmp17_1184 : std_logic_vector(63 downto 0);
    signal tmp18_1189 : std_logic_vector(63 downto 0);
    signal tmp19_1193 : std_logic_vector(31 downto 0);
    signal tmp20_1198 : std_logic_vector(63 downto 0);
    signal tmp21_1204 : std_logic_vector(63 downto 0);
    signal tmp22_1210 : std_logic_vector(0 downto 0);
    signal tmp24_710 : std_logic_vector(31 downto 0);
    signal tmp25_715 : std_logic_vector(31 downto 0);
    signal tmp26_719 : std_logic_vector(31 downto 0);
    signal tmp27_724 : std_logic_vector(31 downto 0);
    signal tmp28_729 : std_logic_vector(63 downto 0);
    signal tmp29_735 : std_logic_vector(63 downto 0);
    signal tmp30_741 : std_logic_vector(0 downto 0);
    signal tmp388_1479 : std_logic_vector(15 downto 0);
    signal tmp389_1603 : std_logic_vector(15 downto 0);
    signal tmp3_1607 : std_logic_vector(31 downto 0);
    signal tmp407_1152 : std_logic_vector(63 downto 0);
    signal tmp408_1158 : std_logic_vector(0 downto 0);
    signal tmp409_1402 : std_logic_vector(63 downto 0);
    signal tmp416_684 : std_logic_vector(31 downto 0);
    signal tmp418_689 : std_logic_vector(31 downto 0);
    signal tmp419_694 : std_logic_vector(63 downto 0);
    signal tmp420_700 : std_logic_vector(63 downto 0);
    signal tmp421_706 : std_logic_vector(0 downto 0);
    signal tmp423_933 : std_logic_vector(63 downto 0);
    signal tmp4_1613 : std_logic_vector(31 downto 0);
    signal tmp6_1617 : std_logic_vector(31 downto 0);
    signal tmp7_1622 : std_logic_vector(15 downto 0);
    signal tmp8_1626 : std_logic_vector(31 downto 0);
    signal tmp9_1631 : std_logic_vector(31 downto 0);
    signal tmp_1006 : std_logic_vector(15 downto 0);
    signal tobool218_1433 : std_logic_vector(0 downto 0);
    signal tobool_964 : std_logic_vector(0 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1010_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1028_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1050_wire : std_logic_vector(63 downto 0);
    signal type_cast_1055_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1061_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1067_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1122_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1127_wire : std_logic_vector(63 downto 0);
    signal type_cast_1130_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1137_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1150_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1156_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1196_wire : std_logic_vector(63 downto 0);
    signal type_cast_1202_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1208_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1215_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1224_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1226_wire : std_logic_vector(63 downto 0);
    signal type_cast_1245_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1263_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1281_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1299_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1317_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1335_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1375_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1400_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1405_wire : std_logic_vector(63 downto 0);
    signal type_cast_1408_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1417_wire : std_logic_vector(63 downto 0);
    signal type_cast_1420_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1425_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1431_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1444_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1454_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1463_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1465_wire : std_logic_vector(15 downto 0);
    signal type_cast_1470_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire : std_logic_vector(63 downto 0);
    signal type_cast_1477_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1523_wire : std_logic_vector(63 downto 0);
    signal type_cast_1528_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1534_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1540_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1580_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1584_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1589_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1595_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1601_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1637_wire : std_logic_vector(31 downto 0);
    signal type_cast_1640_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1673_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1690_wire : std_logic_vector(63 downto 0);
    signal type_cast_1698_wire : std_logic_vector(63 downto 0);
    signal type_cast_1713_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1723_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1733_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1743_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1753_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1763_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_453_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_503_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_528_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_553_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_578_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_603_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_628_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_664_wire : std_logic_vector(63 downto 0);
    signal type_cast_670_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_692_wire : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_704_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_727_wire : std_logic_vector(63 downto 0);
    signal type_cast_733_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_739_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_754_wire : std_logic_vector(63 downto 0);
    signal type_cast_757_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_776_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_794_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_812_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_830_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_848_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_866_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_884_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_931_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_936_wire : std_logic_vector(63 downto 0);
    signal type_cast_939_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_948_wire : std_logic_vector(63 downto 0);
    signal type_cast_951_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_962_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_975_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_981_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_990_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_992_wire : std_logic_vector(15 downto 0);
    signal type_cast_997_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_999_wire : std_logic_vector(63 downto 0);
    signal umax23_1217 : std_logic_vector(63 downto 0);
    signal umax31_748 : std_logic_vector(63 downto 0);
    signal umax422_927 : std_logic_vector(63 downto 0);
    signal umax_1396 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1079_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1079_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1079_resized_base_address <= "00000000000000";
    array_obj_ref_1232_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1232_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1232_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1232_resized_base_address <= "00000000000000";
    array_obj_ref_1552_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1552_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1552_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1552_resized_base_address <= "00000000000000";
    array_obj_ref_763_constant_part_of_offset <= "00000000000000";
    array_obj_ref_763_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_763_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_763_resized_base_address <= "00000000000000";
    ptr_deref_1083_word_offset_0 <= "00000000000000";
    ptr_deref_1369_word_offset_0 <= "00000000000000";
    ptr_deref_1556_word_offset_0 <= "00000000000000";
    ptr_deref_900_word_offset_0 <= "00000000000000";
    type_cast_1004_wire_constant <= "0000000000000001";
    type_cast_1010_wire_constant <= "0000000000000001";
    type_cast_1028_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1055_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1061_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1067_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1122_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1130_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1137_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1150_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1156_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1202_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_1208_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1215_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1224_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1245_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1263_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1281_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1299_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1317_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1335_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1353_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1375_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1400_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1408_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1420_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1425_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1431_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1444_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1454_wire_constant <= "00000000000000000000000000000110";
    type_cast_1463_wire_constant <= "0000000000000000";
    type_cast_1470_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1477_wire_constant <= "0000000000000001";
    type_cast_1483_wire_constant <= "0000000000000001";
    type_cast_1501_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1528_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    type_cast_1534_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1540_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1580_wire_constant <= "11001000";
    type_cast_1584_wire_constant <= "11001000";
    type_cast_1589_wire_constant <= "1111111111111111";
    type_cast_1595_wire_constant <= "1111111111111111";
    type_cast_1601_wire_constant <= "1111111111111111";
    type_cast_1611_wire_constant <= "00000000000000000000000000000001";
    type_cast_1640_wire_constant <= "00000000000000000000000000000000";
    type_cast_1673_wire_constant <= "00000000000000000000000000000001";
    type_cast_1713_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1723_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1733_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1743_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1753_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1763_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1773_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_453_wire_constant <= "00000000000000000000000000001000";
    type_cast_478_wire_constant <= "0000000000001000";
    type_cast_503_wire_constant <= "0000000000001000";
    type_cast_528_wire_constant <= "0000000000001000";
    type_cast_553_wire_constant <= "0000000000001000";
    type_cast_578_wire_constant <= "0000000000001000";
    type_cast_603_wire_constant <= "0000000000001000";
    type_cast_628_wire_constant <= "0000000000001000";
    type_cast_670_wire_constant <= "00000000000000000000000000000011";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_704_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_733_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_739_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_746_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_757_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_776_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_794_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_812_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_830_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_848_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_866_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_884_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_925_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_931_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_939_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_951_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_956_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_962_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_975_wire_constant <= "00000000000000000000000000000001";
    type_cast_981_wire_constant <= "00000000000000000000000000000110";
    type_cast_990_wire_constant <= "0000000000000000";
    type_cast_997_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_1047: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1050_wire;
      req(0) <= phi_stmt_1047_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1047",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1047_ack_0,
          idata => idata,
          odata => shl8x_xix_xlcssa_1047,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1047
    phi_stmt_1220: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1224_wire_constant & type_cast_1226_wire;
      req <= phi_stmt_1220_req_0 & phi_stmt_1220_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1220",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1220_ack_0,
          idata => idata,
          odata => indvar412_1220,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1220
    phi_stmt_1414: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1417_wire & type_cast_1420_wire_constant;
      req <= phi_stmt_1414_req_0 & phi_stmt_1414_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1414",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1414_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1414,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1414
    phi_stmt_1459: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1463_wire_constant & type_cast_1465_wire;
      req <= phi_stmt_1459_req_0 & phi_stmt_1459_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1459",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1459_ack_0,
          idata => idata,
          odata => nx_x022x_xi357_1459,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1459
    phi_stmt_1466: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1470_wire_constant & type_cast_1472_wire;
      req <= phi_stmt_1466_req_0 & phi_stmt_1466_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1466",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1466_ack_0,
          idata => idata,
          odata => elementx_x021x_xi358_1466,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1466
    phi_stmt_1520: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1523_wire;
      req(0) <= phi_stmt_1520_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1520",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1520_ack_0,
          idata => idata,
          odata => shl8x_xi362x_xlcssa_1520,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1520
    phi_stmt_1634: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1637_wire & type_cast_1640_wire_constant;
      req <= phi_stmt_1634_req_0 & phi_stmt_1634_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1634",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1634_ack_0,
          idata => idata,
          odata => indvar_1634,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1634
    phi_stmt_751: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_754_wire & type_cast_757_wire_constant;
      req <= phi_stmt_751_req_0 & phi_stmt_751_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_751",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_751_ack_0,
          idata => idata,
          odata => indvar426_751,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_751
    phi_stmt_945: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_948_wire & type_cast_951_wire_constant;
      req <= phi_stmt_945_req_0 & phi_stmt_945_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_945",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_945_ack_0,
          idata => idata,
          odata => ix_x0x_xlcssa_945,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_945
    phi_stmt_986: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_990_wire_constant & type_cast_992_wire;
      req <= phi_stmt_986_req_0 & phi_stmt_986_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_986",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_986_ack_0,
          idata => idata,
          odata => nx_x022x_xi_986,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_986
    phi_stmt_993: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_997_wire_constant & type_cast_999_wire;
      req <= phi_stmt_993_req_0 & phi_stmt_993_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_993",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_993_ack_0,
          idata => idata,
          odata => elementx_x021x_xi_993,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_993
    -- flow-through select operator MUX_1216_inst
    umax23_1217 <= tmp21_1204 when (tmp22_1210(0) /=  '0') else type_cast_1215_wire_constant;
    -- flow-through select operator MUX_1395_inst
    umax_1396 <= tmp407_1152 when (tmp408_1158(0) /=  '0') else type_cast_1394_wire_constant;
    -- flow-through select operator MUX_747_inst
    umax31_748 <= tmp29_735 when (tmp30_741(0) /=  '0') else type_cast_746_wire_constant;
    -- flow-through select operator MUX_926_inst
    umax422_927 <= tmp420_700 when (tmp421_706(0) /=  '0') else type_cast_925_wire_constant;
    addr_of_1080_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1080_final_reg_req_0;
      addr_of_1080_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1080_final_reg_req_1;
      addr_of_1080_final_reg_ack_1<= rack(0);
      addr_of_1080_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1080_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1079_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx143_1081,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1233_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1233_final_reg_req_0;
      addr_of_1233_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1233_final_reg_req_1;
      addr_of_1233_final_reg_ack_1<= rack(0);
      addr_of_1233_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1233_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1232_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1234,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1553_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1553_final_reg_req_0;
      addr_of_1553_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1553_final_reg_req_1;
      addr_of_1553_final_reg_ack_1<= rack(0);
      addr_of_1553_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1553_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1552_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx226_1554,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_764_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_764_final_reg_req_0;
      addr_of_764_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_764_final_reg_req_1;
      addr_of_764_final_reg_ack_1<= rack(0);
      addr_of_764_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_764_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_763_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1018_inst_req_0;
      type_cast_1018_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1018_inst_req_1;
      type_cast_1018_inst_ack_1<= rack(0);
      type_cast_1018_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1015,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1033_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1033_inst_req_0;
      type_cast_1033_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1033_inst_req_1;
      type_cast_1033_inst_ack_1<= rack(0);
      type_cast_1033_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1033_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1006,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi_1034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1050_inst_req_0;
      type_cast_1050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1050_inst_req_1;
      type_cast_1050_inst_ack_1<= rack(0);
      type_cast_1050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1050_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1090_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1090_inst_req_0;
      type_cast_1090_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1090_inst_req_1;
      type_cast_1090_inst_ack_1<= rack(0);
      type_cast_1090_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1090_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv145_1091,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1094_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1094_inst_req_0;
      type_cast_1094_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1094_inst_req_1;
      type_cast_1094_inst_ack_1<= rack(0);
      type_cast_1094_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1094_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_1095,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1098_inst_req_0;
      type_cast_1098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1098_inst_req_1;
      type_cast_1098_inst_ack_1<= rack(0);
      type_cast_1098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv150_1099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1102_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1102_inst_req_0;
      type_cast_1102_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1102_inst_req_1;
      type_cast_1102_inst_ack_1<= rack(0);
      type_cast_1102_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1102_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1127_inst
    process(sext_1124) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := sext_1124(63 downto 0);
      type_cast_1127_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1132_inst
    process(ASHR_i64_i64_1131_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1131_wire(63 downto 0);
      conv155_1133 <= tmp_var; -- 
    end process;
    type_cast_1161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1161_inst_req_0;
      type_cast_1161_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1161_inst_req_1;
      type_cast_1161_inst_ack_1<= rack(0);
      type_cast_1161_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_592,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1162,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1165_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1165_inst_req_0;
      type_cast_1165_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1165_inst_req_1;
      type_cast_1165_inst_ack_1<= rack(0);
      type_cast_1165_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1165_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp13_1166,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1174_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1174_inst_req_0;
      type_cast_1174_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1174_inst_req_1;
      type_cast_1174_inst_ack_1<= rack(0);
      type_cast_1174_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1174_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_1175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1183_inst_req_0;
      type_cast_1183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1183_inst_req_1;
      type_cast_1183_inst_ack_1<= rack(0);
      type_cast_1183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_642,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp17_1184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1192_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1192_inst_req_0;
      type_cast_1192_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1192_inst_req_1;
      type_cast_1192_inst_ack_1<= rack(0);
      type_cast_1192_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1192_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp18_1189,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp19_1193,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1197_inst_req_0;
      type_cast_1197_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1197_inst_req_1;
      type_cast_1197_inst_ack_1<= rack(0);
      type_cast_1197_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1196_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1198,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1226_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1226_inst_req_0;
      type_cast_1226_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1226_inst_req_1;
      type_cast_1226_inst_ack_1<= rack(0);
      type_cast_1226_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1226_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext413_1377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1226_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1240_inst_req_0;
      type_cast_1240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1240_inst_req_1;
      type_cast_1240_inst_ack_1<= rack(0);
      type_cast_1240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call164_1237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_1241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1253_inst_req_0;
      type_cast_1253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1253_inst_req_1;
      type_cast_1253_inst_ack_1<= rack(0);
      type_cast_1253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1271_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1271_inst_req_0;
      type_cast_1271_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1271_inst_req_1;
      type_cast_1271_inst_ack_1<= rack(0);
      type_cast_1271_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1271_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1268,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1272,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1289_inst_req_0;
      type_cast_1289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1289_inst_req_1;
      type_cast_1289_inst_ack_1<= rack(0);
      type_cast_1289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1290,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1307_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1307_inst_req_0;
      type_cast_1307_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1307_inst_req_1;
      type_cast_1307_inst_ack_1<= rack(0);
      type_cast_1307_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1307_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1304,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1308,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1325_inst_req_0;
      type_cast_1325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1325_inst_req_1;
      type_cast_1325_inst_ack_1<= rack(0);
      type_cast_1325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1325_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1322,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1326,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1343_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1343_inst_req_0;
      type_cast_1343_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1343_inst_req_1;
      type_cast_1343_inst_ack_1<= rack(0);
      type_cast_1343_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1343_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call198_1340,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv200_1344,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1361_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1361_inst_req_0;
      type_cast_1361_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1361_inst_req_1;
      type_cast_1361_inst_ack_1<= rack(0);
      type_cast_1361_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1361_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call204_1358,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv206_1362,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1405_inst
    process(tmp409_1402) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp409_1402(63 downto 0);
      type_cast_1405_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1410_inst
    process(ASHR_i64_i64_1409_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_1409_wire(63 downto 0);
      phitmp387_1411 <= tmp_var; -- 
    end process;
    type_cast_1417_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1417_inst_req_0;
      type_cast_1417_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1417_inst_req_1;
      type_cast_1417_inst_ack_1<= rack(0);
      type_cast_1417_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1417_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp387_1411,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1417_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1449_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1449_inst_req_0;
      type_cast_1449_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1449_inst_req_1;
      type_cast_1449_inst_ack_1<= rack(0);
      type_cast_1449_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1449_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_57_1446,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv2x_xi354_1450,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1465_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1465_inst_req_0;
      type_cast_1465_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1465_inst_req_1;
      type_cast_1465_inst_ack_1<= rack(0);
      type_cast_1465_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1465_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_65_1485,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1465_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1472_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1472_inst_req_0;
      type_cast_1472_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1472_inst_req_1;
      type_cast_1472_inst_ack_1<= rack(0);
      type_cast_1472_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1472_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_1503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1472_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1491_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1491_inst_req_0;
      type_cast_1491_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1491_inst_req_1;
      type_cast_1491_inst_ack_1<= rack(0);
      type_cast_1491_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1491_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi359_1488,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi360_1492,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1506_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1506_inst_req_0;
      type_cast_1506_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1506_inst_req_1;
      type_cast_1506_inst_ack_1<= rack(0);
      type_cast_1506_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1506_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp388_1479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => convx_xi363_1507,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1523_inst_req_0;
      type_cast_1523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1523_inst_req_1;
      type_cast_1523_inst_ack_1<= rack(0);
      type_cast_1523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi362_1503,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1523_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1606_inst_req_0;
      type_cast_1606_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1606_inst_req_1;
      type_cast_1606_inst_ack_1<= rack(0);
      type_cast_1606_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1606_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp389_1603,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1616_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1616_inst_req_0;
      type_cast_1616_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1616_inst_req_1;
      type_cast_1616_inst_ack_1<= rack(0);
      type_cast_1616_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1616_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add63_617,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp6_1617,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1625_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1625_inst_req_0;
      type_cast_1625_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1625_inst_req_1;
      type_cast_1625_inst_ack_1<= rack(0);
      type_cast_1625_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1625_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp7_1622,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp8_1626,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1637_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1637_inst_req_0;
      type_cast_1637_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1637_inst_req_1;
      type_cast_1637_inst_ack_1<= rack(0);
      type_cast_1637_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1637_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1675,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1637_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1654_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1654_inst_req_0;
      type_cast_1654_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1654_inst_req_1;
      type_cast_1654_inst_ack_1<= rack(0);
      type_cast_1654_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1654_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul254_1646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv255_1655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1658_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1658_inst_req_0;
      type_cast_1658_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1658_inst_req_1;
      type_cast_1658_inst_ack_1<= rack(0);
      type_cast_1658_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1658_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul260_1651,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv261_1659,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1691_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1691_inst_req_0;
      type_cast_1691_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1691_inst_req_1;
      type_cast_1691_inst_ack_1<= rack(0);
      type_cast_1691_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1691_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1690_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv230_1692,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1699_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1699_inst_req_0;
      type_cast_1699_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1699_inst_req_1;
      type_cast_1699_inst_ack_1<= rack(0);
      type_cast_1699_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1699_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1698_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv285_1700,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1708_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1708_inst_req_0;
      type_cast_1708_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1708_inst_req_1;
      type_cast_1708_inst_ack_1<= rack(0);
      type_cast_1708_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1708_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub289_1705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv293_1709,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1718_inst_req_0;
      type_cast_1718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1718_inst_req_1;
      type_cast_1718_inst_ack_1<= rack(0);
      type_cast_1718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr296_1715,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv299_1719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1728_inst_req_0;
      type_cast_1728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1728_inst_req_1;
      type_cast_1728_inst_ack_1<= rack(0);
      type_cast_1728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr302_1725,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv305_1729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1738_inst_req_0;
      type_cast_1738_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1738_inst_req_1;
      type_cast_1738_inst_ack_1<= rack(0);
      type_cast_1738_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1738_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr308_1735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv311_1739,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1748_inst_req_0;
      type_cast_1748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1748_inst_req_1;
      type_cast_1748_inst_ack_1<= rack(0);
      type_cast_1748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr314_1745,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv317_1749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1758_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1758_inst_req_0;
      type_cast_1758_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1758_inst_req_1;
      type_cast_1758_inst_ack_1<= rack(0);
      type_cast_1758_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1758_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr320_1755,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv323_1759,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1768_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1768_inst_req_0;
      type_cast_1768_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1768_inst_req_1;
      type_cast_1768_inst_ack_1<= rack(0);
      type_cast_1768_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1768_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr326_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv329_1769,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1778_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1778_inst_req_0;
      type_cast_1778_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1778_inst_req_1;
      type_cast_1778_inst_ack_1<= rack(0);
      type_cast_1778_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1778_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr332_1775,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv335_1779,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_448_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_448_inst_req_0;
      type_cast_448_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_448_inst_req_1;
      type_cast_448_inst_ack_1<= rack(0);
      type_cast_448_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_448_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_445,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_449,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_461_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_461_inst_req_0;
      type_cast_461_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_461_inst_req_1;
      type_cast_461_inst_ack_1<= rack(0);
      type_cast_461_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_461_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_458,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_462,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_473_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_473_inst_req_0;
      type_cast_473_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_473_inst_req_1;
      type_cast_473_inst_ack_1<= rack(0);
      type_cast_473_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_473_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_470,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_474,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_498_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_498_inst_req_0;
      type_cast_498_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_498_inst_req_1;
      type_cast_498_inst_ack_1<= rack(0);
      type_cast_498_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_498_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_495,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_499,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_511_inst_req_0;
      type_cast_511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_511_inst_req_1;
      type_cast_511_inst_ack_1<= rack(0);
      type_cast_511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_508,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_523_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_523_inst_req_0;
      type_cast_523_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_523_inst_req_1;
      type_cast_523_inst_ack_1<= rack(0);
      type_cast_523_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_523_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_520,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_524,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_536_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_536_inst_req_0;
      type_cast_536_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_536_inst_req_1;
      type_cast_536_inst_ack_1<= rack(0);
      type_cast_536_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_536_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_533,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_537,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_548_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_548_inst_req_0;
      type_cast_548_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_548_inst_req_1;
      type_cast_548_inst_ack_1<= rack(0);
      type_cast_548_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_548_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_545,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_549,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_573_inst_req_0;
      type_cast_573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_573_inst_req_1;
      type_cast_573_inst_ack_1<= rack(0);
      type_cast_573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_570,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_586_inst_req_0;
      type_cast_586_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_586_inst_req_1;
      type_cast_586_inst_ack_1<= rack(0);
      type_cast_586_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_586_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_583,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_587,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_598_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_598_inst_req_0;
      type_cast_598_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_598_inst_req_1;
      type_cast_598_inst_ack_1<= rack(0);
      type_cast_598_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_598_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_595,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_599,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_611_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_611_inst_req_0;
      type_cast_611_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_611_inst_req_1;
      type_cast_611_inst_ack_1<= rack(0);
      type_cast_611_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_611_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_608,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_612,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_623_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_623_inst_req_0;
      type_cast_623_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_623_inst_req_1;
      type_cast_623_inst_ack_1<= rack(0);
      type_cast_623_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_623_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_620,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_624,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_636_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_636_inst_req_1;
      type_cast_636_inst_ack_1<= rack(0);
      type_cast_636_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_636_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_633,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_637,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_645_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_645_inst_req_0;
      type_cast_645_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_645_inst_req_1;
      type_cast_645_inst_ack_1<= rack(0);
      type_cast_645_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_645_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_646,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_665_inst_req_0;
      type_cast_665_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_665_inst_req_1;
      type_cast_665_inst_ack_1<= rack(0);
      type_cast_665_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_665_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_664_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv83_666,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_693_inst_req_0;
      type_cast_693_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_693_inst_req_1;
      type_cast_693_inst_ack_1<= rack(0);
      type_cast_693_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_693_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_692_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp419_694,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_709_inst_req_0;
      type_cast_709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_709_inst_req_1;
      type_cast_709_inst_ack_1<= rack(0);
      type_cast_709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp24_710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_718_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_718_inst_req_0;
      type_cast_718_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_718_inst_req_1;
      type_cast_718_inst_ack_1<= rack(0);
      type_cast_718_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_718_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_517,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp26_719,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_728_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_728_inst_req_0;
      type_cast_728_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_728_inst_req_1;
      type_cast_728_inst_ack_1<= rack(0);
      type_cast_728_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_728_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_727_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp28_729,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_754_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_754_inst_req_0;
      type_cast_754_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_754_inst_req_1;
      type_cast_754_inst_ack_1<= rack(0);
      type_cast_754_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_754_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext427_908,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_754_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_771_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_771_inst_req_0;
      type_cast_771_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_771_inst_req_1;
      type_cast_771_inst_ack_1<= rack(0);
      type_cast_771_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_771_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_768,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_772,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_784_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_784_inst_req_0;
      type_cast_784_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_784_inst_req_1;
      type_cast_784_inst_ack_1<= rack(0);
      type_cast_784_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_784_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call93_781,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv95_785,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_802_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_802_inst_req_0;
      type_cast_802_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_802_inst_req_1;
      type_cast_802_inst_ack_1<= rack(0);
      type_cast_802_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_802_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call99_799,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv101_803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_820_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_820_inst_req_0;
      type_cast_820_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_820_inst_req_1;
      type_cast_820_inst_ack_1<= rack(0);
      type_cast_820_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_820_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call105_817,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv107_821,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_838_inst_req_0;
      type_cast_838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_838_inst_req_1;
      type_cast_838_inst_ack_1<= rack(0);
      type_cast_838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call111_835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv113_839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_856_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_856_inst_req_0;
      type_cast_856_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_856_inst_req_1;
      type_cast_856_inst_ack_1<= rack(0);
      type_cast_856_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_856_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call117_853,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv119_857,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_874_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_874_inst_req_0;
      type_cast_874_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_874_inst_req_1;
      type_cast_874_inst_ack_1<= rack(0);
      type_cast_874_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_874_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call123_871,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv125_875,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_892_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_892_inst_req_0;
      type_cast_892_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_892_inst_req_1;
      type_cast_892_inst_ack_1<= rack(0);
      type_cast_892_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_892_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_889,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv131_893,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_936_inst
    process(tmp423_933) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := tmp423_933(63 downto 0);
      type_cast_936_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_941_inst
    process(ASHR_i64_i64_940_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := ASHR_i64_i64_940_wire(63 downto 0);
      phitmp_942 <= tmp_var; -- 
    end process;
    type_cast_948_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_948_inst_req_0;
      type_cast_948_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_948_inst_req_1;
      type_cast_948_inst_ack_1<= rack(0);
      type_cast_948_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_948_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp_942,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_948_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_992_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_992_inst_req_0;
      type_cast_992_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_992_inst_req_1;
      type_cast_992_inst_ack_1<= rack(0);
      type_cast_992_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_992_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => iNsTr_35_1012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_992_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_999_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_999_inst_req_0;
      type_cast_999_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_999_inst_req_1;
      type_cast_999_inst_ack_1<= rack(0);
      type_cast_999_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_999_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shl8x_xi_1030,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_999_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1079_index_1_rename
    process(R_ix_x0x_xlcssa_1078_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x0x_xlcssa_1078_resized;
      ov(13 downto 0) := iv;
      R_ix_x0x_xlcssa_1078_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_index_1_resize
    process(ix_x0x_xlcssa_945) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x0x_xlcssa_945;
      ov := iv(13 downto 0);
      R_ix_x0x_xlcssa_1078_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1079_root_address_inst
    process(array_obj_ref_1079_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1079_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1079_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1232_index_1_rename
    process(R_indvar412_1231_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar412_1231_resized;
      ov(13 downto 0) := iv;
      R_indvar412_1231_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1232_index_1_resize
    process(indvar412_1220) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar412_1220;
      ov := iv(13 downto 0);
      R_indvar412_1231_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1232_root_address_inst
    process(array_obj_ref_1232_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1232_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1232_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1552_index_1_rename
    process(R_ix_x1x_xlcssa_1551_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1551_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1551_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1552_index_1_resize
    process(ix_x1x_xlcssa_1414) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1414;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1551_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1552_root_address_inst
    process(array_obj_ref_1552_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1552_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1552_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_763_index_1_rename
    process(R_indvar426_762_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar426_762_resized;
      ov(13 downto 0) := iv;
      R_indvar426_762_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_763_index_1_resize
    process(indvar426_751) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar426_751;
      ov := iv(13 downto 0);
      R_indvar426_762_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_763_root_address_inst
    process(array_obj_ref_763_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_763_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_763_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1083_addr_0
    process(ptr_deref_1083_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1083_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1083_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1083_base_resize
    process(arrayidx143_1081) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx143_1081;
      ov := iv(13 downto 0);
      ptr_deref_1083_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1083_gather_scatter
    process(shl14x_xi_1074) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi_1074;
      ov(63 downto 0) := iv;
      ptr_deref_1083_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1083_root_address_inst
    process(ptr_deref_1083_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1083_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1083_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1369_addr_0
    process(ptr_deref_1369_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1369_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1369_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1369_base_resize
    process(arrayidx211_1234) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1234;
      ov := iv(13 downto 0);
      ptr_deref_1369_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1369_gather_scatter
    process(add207_1367) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add207_1367;
      ov(63 downto 0) := iv;
      ptr_deref_1369_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1369_root_address_inst
    process(ptr_deref_1369_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1369_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1369_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1556_addr_0
    process(ptr_deref_1556_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1556_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1556_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1556_base_resize
    process(arrayidx226_1554) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx226_1554;
      ov := iv(13 downto 0);
      ptr_deref_1556_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1556_gather_scatter
    process(shl14x_xi372_1547) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl14x_xi372_1547;
      ov(63 downto 0) := iv;
      ptr_deref_1556_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1556_root_address_inst
    process(ptr_deref_1556_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1556_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1556_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_900_addr_0
    process(ptr_deref_900_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_900_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_900_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_900_base_resize
    process(arrayidx_765) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_765;
      ov := iv(13 downto 0);
      ptr_deref_900_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_900_gather_scatter
    process(add132_898) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add132_898;
      ov(63 downto 0) := iv;
      ptr_deref_900_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_900_root_address_inst
    process(ptr_deref_900_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_900_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_900_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1040_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi_1039;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1040_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1040_branch_req_0,
          ack0 => if_stmt_1040_branch_ack_0,
          ack1 => if_stmt_1040_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1140_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp161379_1139;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1140_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1140_branch_req_0,
          ack0 => if_stmt_1140_branch_ack_0,
          ack1 => if_stmt_1140_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1383_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1382;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1383_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1383_branch_req_0,
          ack0 => if_stmt_1383_branch_ack_0,
          ack1 => if_stmt_1383_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1434_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool218_1433;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1434_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1434_branch_req_0,
          ack0 => if_stmt_1434_branch_ack_0,
          ack1 => if_stmt_1434_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1513_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmpx_xi364_1512;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1513_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1513_branch_req_0,
          ack0 => if_stmt_1513_branch_ack_0,
          ack1 => if_stmt_1513_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1681_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond5_1680;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1681_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1681_branch_req_0,
          ack0 => if_stmt_1681_branch_ack_0,
          ack1 => if_stmt_1681_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_673_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp383_672;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_673_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_673_branch_req_0,
          ack0 => if_stmt_673_branch_ack_0,
          ack1 => if_stmt_673_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_914_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond32_913;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_914_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_914_branch_req_0,
          ack0 => if_stmt_914_branch_ack_0,
          ack1 => if_stmt_914_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_965_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_964;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_965_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_965_branch_req_0,
          ack0 => if_stmt_965_branch_ack_0,
          ack1 => if_stmt_965_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1005_inst
    process(nx_x022x_xi_986) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_986, type_cast_1004_wire_constant, tmp_var);
      tmp_1006 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1011_inst
    process(nx_x022x_xi_986) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi_986, type_cast_1010_wire_constant, tmp_var);
      iNsTr_35_1012 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1478_inst
    process(nx_x022x_xi357_1459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_1459, type_cast_1477_wire_constant, tmp_var);
      tmp388_1479 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1484_inst
    process(nx_x022x_xi357_1459) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x022x_xi357_1459, type_cast_1483_wire_constant, tmp_var);
      iNsTr_65_1485 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1590_inst
    process(add43_567) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add43_567, type_cast_1589_wire_constant, tmp_var);
      sub_1591 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1596_inst
    process(add63_617) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add63_617, type_cast_1595_wire_constant, tmp_var);
      sub269_1597 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1602_inst
    process(add53_592) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_592, type_cast_1601_wire_constant, tmp_var);
      tmp389_1603 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1612_inst
    process(tmp3_1607) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1607, type_cast_1611_wire_constant, tmp_var);
      tmp4_1613 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1650_inst
    process(tmp9_1631, mul254_1646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp9_1631, mul254_1646, tmp_var);
      mul260_1651 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1674_inst
    process(indvar_1634) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1634, type_cast_1673_wire_constant, tmp_var);
      indvarx_xnext_1675 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1376_inst
    process(indvar412_1220) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar412_1220, type_cast_1375_wire_constant, tmp_var);
      indvarx_xnext413_1377 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_907_inst
    process(indvar426_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar426_751, type_cast_906_wire_constant, tmp_var);
      indvarx_xnext427_908 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1455_inst
    process(conv2x_xi354_1450) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi354_1450, type_cast_1454_wire_constant, tmp_var);
      shlx_xi355_1456 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_982_inst
    process(conv2x_xi_977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv2x_xi_977, type_cast_981_wire_constant, tmp_var);
      shlx_xi_983 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1062_inst
    process(Bx_xnot_1057) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(Bx_xnot_1057, type_cast_1061_wire_constant, tmp_var);
      add1216x_xi_1063 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1426_inst
    process(conv155_1133) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv155_1133, type_cast_1425_wire_constant, tmp_var);
      and217_1427 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1535_inst
    process(iNsTr_87_1530) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(iNsTr_87_1530, type_cast_1534_wire_constant, tmp_var);
      add1216x_xi370_1536 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_957_inst
    process(conv83_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv83_666, type_cast_956_wire_constant, tmp_var);
      and_958 <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1131_inst
    process(type_cast_1127_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1127_wire, type_cast_1130_wire_constant, tmp_var);
      ASHR_i64_i64_1131_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_1409_inst
    process(type_cast_1405_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1405_wire, type_cast_1408_wire_constant, tmp_var);
      ASHR_i64_i64_1409_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i64_i64_940_inst
    process(type_cast_936_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_936_wire, type_cast_939_wire_constant, tmp_var);
      ASHR_i64_i64_940_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1679_inst
    process(indvarx_xnext_1675, tmp4_1613) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1675, tmp4_1613, tmp_var);
      exitcond5_1680 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1381_inst
    process(indvarx_xnext413_1377, umax23_1217) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext413_1377, umax23_1217, tmp_var);
      exitcond_1382 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1432_inst
    process(and217_1427) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and217_1427, type_cast_1431_wire_constant, tmp_var);
      tobool218_1433 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_912_inst
    process(indvarx_xnext427_908, umax31_748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext427_908, umax31_748, tmp_var);
      exitcond32_913 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_963_inst
    process(and_958) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_958, type_cast_962_wire_constant, tmp_var);
      tobool_964 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1151_inst
    process(conv155_1133) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(conv155_1133, type_cast_1150_wire_constant, tmp_var);
      tmp407_1152 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1203_inst
    process(tmp20_1198) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp20_1198, type_cast_1202_wire_constant, tmp_var);
      tmp21_1204 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1714_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1713_wire_constant, tmp_var);
      shr296_1715 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1724_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1723_wire_constant, tmp_var);
      shr302_1725 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1734_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1733_wire_constant, tmp_var);
      shr308_1735 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1744_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1743_wire_constant, tmp_var);
      shr314_1745 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1754_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1753_wire_constant, tmp_var);
      shr320_1755 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1764_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1763_wire_constant, tmp_var);
      shr326_1765 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1774_inst
    process(sub289_1705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub289_1705, type_cast_1773_wire_constant, tmp_var);
      shr332_1775 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_699_inst
    process(tmp419_694) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp419_694, type_cast_698_wire_constant, tmp_var);
      tmp420_700 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_734_inst
    process(tmp28_729) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp28_729, type_cast_733_wire_constant, tmp_var);
      tmp29_735 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1568_inst
    process(add73_642, add23_517) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_642, add23_517, tmp_var);
      mul236_1569 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1573_inst
    process(add43_567, add33_542) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add43_567, add33_542, tmp_var);
      mul249_1574 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1621_inst
    process(add73_642, add23_517) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_642, add23_517, tmp_var);
      tmp7_1622 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1630_inst
    process(tmp6_1617, tmp8_1626) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp6_1617, tmp8_1626, tmp_var);
      tmp9_1631 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1645_inst
    process(tmp9_1631, indvar_1634) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp9_1631, indvar_1634, tmp_var);
      mul254_1646 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_654_inst
    process(conv79_646, add_467) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_646, add_467, tmp_var);
      mul_655 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_659_inst
    process(mul_655, conv81_650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_655, conv81_650, tmp_var);
      mul82_660 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_683_inst
    process(add_467, conv79_646) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_467, conv79_646, tmp_var);
      tmp416_684 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_688_inst
    process(tmp416_684, conv81_650) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp416_684, conv81_650, tmp_var);
      tmp418_689 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_714_inst
    process(add_467, tmp24_710) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_467, tmp24_710, tmp_var);
      tmp25_715 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_723_inst
    process(tmp25_715, tmp26_719) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp25_715, tmp26_719, tmp_var);
      tmp27_724 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1107_inst
    process(conv153_1103, conv145_1091) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv153_1103, conv145_1091, tmp_var);
      mul148_1108 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1112_inst
    process(mul148_1108, conv150_1099) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul148_1108, conv150_1099, tmp_var);
      mul151_1113 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1117_inst
    process(mul151_1113, conv147_1095) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul151_1113, conv147_1095, tmp_var);
      mul154_1118 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1170_inst
    process(tmp12_1162, tmp13_1166) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_1162, tmp13_1166, tmp_var);
      tmp14_1171 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1179_inst
    process(tmp14_1171, tmp15_1175) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_1171, tmp15_1175, tmp_var);
      tmp16_1180 <= tmp_var; --
    end process;
    -- binary operator MUL_u64_u64_1188_inst
    process(tmp16_1180, tmp17_1184) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp16_1180, tmp17_1184, tmp_var);
      tmp18_1189 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_491_inst
    process(shl10_480, conv12_487) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_480, conv12_487, tmp_var);
      add13_492 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_516_inst
    process(shl20_505, conv22_512) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_505, conv22_512, tmp_var);
      add23_517 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_541_inst
    process(shl30_530, conv32_537) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_530, conv32_537, tmp_var);
      add33_542 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_566_inst
    process(shl40_555, conv42_562) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_555, conv42_562, tmp_var);
      add43_567 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_591_inst
    process(shl50_580, conv52_587) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_580, conv52_587, tmp_var);
      add53_592 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_616_inst
    process(shl60_605, conv62_612) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_605, conv62_612, tmp_var);
      add63_617 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_641_inst
    process(shl70_630, conv72_637) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_630, conv72_637, tmp_var);
      add73_642 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_466_inst
    process(shl_455, conv3_462) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_455, conv3_462, tmp_var);
      add_467 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1023_inst
    process(conv5x_xi_1019, elementx_x021x_xi_993) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1019, elementx_x021x_xi_993, tmp_var);
      addx_xi_1024 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1258_inst
    process(shl167_1247, conv170_1254) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1247, conv170_1254, tmp_var);
      add171_1259 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1276_inst
    process(shl173_1265, conv176_1272) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1265, conv176_1272, tmp_var);
      add177_1277 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1294_inst
    process(shl179_1283, conv182_1290) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1283, conv182_1290, tmp_var);
      add183_1295 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1312_inst
    process(shl185_1301, conv188_1308) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1301, conv188_1308, tmp_var);
      add189_1313 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1330_inst
    process(shl191_1319, conv194_1326) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1319, conv194_1326, tmp_var);
      add195_1331 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1348_inst
    process(shl197_1337, conv200_1344) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl197_1337, conv200_1344, tmp_var);
      add201_1349 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1366_inst
    process(shl203_1355, conv206_1362) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl203_1355, conv206_1362, tmp_var);
      add207_1367 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1496_inst
    process(conv5x_xi360_1492, elementx_x021x_xi358_1466) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi360_1492, elementx_x021x_xi358_1466, tmp_var);
      addx_xi361_1497 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_789_inst
    process(shl92_778, conv95_785) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl92_778, conv95_785, tmp_var);
      add96_790 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_807_inst
    process(shl98_796, conv101_803) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl98_796, conv101_803, tmp_var);
      add102_808 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_825_inst
    process(shl104_814, conv107_821) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl104_814, conv107_821, tmp_var);
      add108_826 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_843_inst
    process(shl110_832, conv113_839) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl110_832, conv113_839, tmp_var);
      add114_844 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_861_inst
    process(shl116_850, conv119_857) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl116_850, conv119_857, tmp_var);
      add120_862 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_879_inst
    process(shl122_868, conv125_875) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl122_868, conv125_875, tmp_var);
      add126_880 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_897_inst
    process(shl128_886, conv131_893) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl128_886, conv131_893, tmp_var);
      add132_898 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_479_inst
    process(conv9_474) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_474, type_cast_478_wire_constant, tmp_var);
      shl10_480 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_504_inst
    process(conv19_499) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_499, type_cast_503_wire_constant, tmp_var);
      shl20_505 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_529_inst
    process(conv29_524) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_524, type_cast_528_wire_constant, tmp_var);
      shl30_530 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_554_inst
    process(conv39_549) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_549, type_cast_553_wire_constant, tmp_var);
      shl40_555 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_579_inst
    process(conv49_574) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_574, type_cast_578_wire_constant, tmp_var);
      shl50_580 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_604_inst
    process(conv59_599) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_599, type_cast_603_wire_constant, tmp_var);
      shl60_605 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_629_inst
    process(conv69_624) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_624, type_cast_628_wire_constant, tmp_var);
      shl70_630 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_454_inst
    process(conv1_449) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_449, type_cast_453_wire_constant, tmp_var);
      shl_455 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_976_inst
    process(mul82_660) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul82_660, type_cast_975_wire_constant, tmp_var);
      conv2x_xi_977 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1029_inst
    process(addx_xi_1024) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1024, type_cast_1028_wire_constant, tmp_var);
      shl8x_xi_1030 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1056_inst
    process(conv83_666) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv83_666, type_cast_1055_wire_constant, tmp_var);
      Bx_xnot_1057 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1073_inst
    process(shl8x_xix_xlcssa_1047, sh_promx_xi_1069) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xix_xlcssa_1047, sh_promx_xi_1069, tmp_var);
      shl14x_xi_1074 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1123_inst
    process(mul154_1118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1118, type_cast_1122_wire_constant, tmp_var);
      sext_1124 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1246_inst
    process(conv165_1241) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv165_1241, type_cast_1245_wire_constant, tmp_var);
      shl167_1247 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1264_inst
    process(add171_1259) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1259, type_cast_1263_wire_constant, tmp_var);
      shl173_1265 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1282_inst
    process(add177_1277) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1277, type_cast_1281_wire_constant, tmp_var);
      shl179_1283 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1300_inst
    process(add183_1295) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1295, type_cast_1299_wire_constant, tmp_var);
      shl185_1301 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1318_inst
    process(add189_1313) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1313, type_cast_1317_wire_constant, tmp_var);
      shl191_1319 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1336_inst
    process(add195_1331) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add195_1331, type_cast_1335_wire_constant, tmp_var);
      shl197_1337 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1354_inst
    process(add201_1349) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add201_1349, type_cast_1353_wire_constant, tmp_var);
      shl203_1355 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1401_inst
    process(umax_1396) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax_1396, type_cast_1400_wire_constant, tmp_var);
      tmp409_1402 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1445_inst
    process(mul154_1118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1118, type_cast_1444_wire_constant, tmp_var);
      iNsTr_57_1446 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1502_inst
    process(addx_xi361_1497) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi361_1497, type_cast_1501_wire_constant, tmp_var);
      shl8x_xi362_1503 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1529_inst
    process(mul154_1118) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(mul154_1118, type_cast_1528_wire_constant, tmp_var);
      iNsTr_87_1530 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1546_inst
    process(shl8x_xi362x_xlcssa_1520, sh_promx_xi371_1542) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shl8x_xi362x_xlcssa_1520, sh_promx_xi371_1542, tmp_var);
      shl14x_xi372_1547 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_777_inst
    process(conv90_772) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv90_772, type_cast_776_wire_constant, tmp_var);
      shl92_778 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_795_inst
    process(add96_790) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add96_790, type_cast_794_wire_constant, tmp_var);
      shl98_796 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_813_inst
    process(add102_808) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add102_808, type_cast_812_wire_constant, tmp_var);
      shl104_814 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_831_inst
    process(add108_826) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add108_826, type_cast_830_wire_constant, tmp_var);
      shl110_832 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_849_inst
    process(add114_844) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add114_844, type_cast_848_wire_constant, tmp_var);
      shl116_850 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_867_inst
    process(add120_862) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add120_862, type_cast_866_wire_constant, tmp_var);
      shl122_868 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_885_inst
    process(add126_880) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add126_880, type_cast_884_wire_constant, tmp_var);
      shl128_886 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_932_inst
    process(umax422_927) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(umax422_927, type_cast_931_wire_constant, tmp_var);
      tmp423_933 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1704_inst
    process(conv285_1700, conv230_1692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv285_1700, conv230_1692, tmp_var);
      sub289_1705 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_671_inst
    process(mul82_660) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_660, type_cast_670_wire_constant, tmp_var);
      cmp383_672 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1138_inst
    process(conv155_1133) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(conv155_1133, type_cast_1137_wire_constant, tmp_var);
      cmp161379_1139 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1157_inst
    process(tmp407_1152) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp407_1152, type_cast_1156_wire_constant, tmp_var);
      tmp408_1158 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_1209_inst
    process(tmp21_1204) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp21_1204, type_cast_1208_wire_constant, tmp_var);
      tmp22_1210 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_705_inst
    process(tmp420_700) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp420_700, type_cast_704_wire_constant, tmp_var);
      tmp421_706 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_740_inst
    process(tmp29_735) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp29_735, type_cast_739_wire_constant, tmp_var);
      tmp30_741 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1038_inst
    process(convx_xi_1034, shlx_xi_983) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi_1034, shlx_xi_983, tmp_var);
      cmpx_xi_1039 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1511_inst
    process(convx_xi363_1507, shlx_xi355_1456) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(convx_xi363_1507, shlx_xi355_1456, tmp_var);
      cmpx_xi364_1512 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1068_inst
    process(add1216x_xi_1063) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi_1063, type_cast_1067_wire_constant, tmp_var);
      sh_promx_xi_1069 <= tmp_var; --
    end process;
    -- binary operator XOR_u64_u64_1541_inst
    process(add1216x_xi370_1536) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntXor_proc(add1216x_xi370_1536, type_cast_1540_wire_constant, tmp_var);
      sh_promx_xi371_1542 <= tmp_var; --
    end process;
    -- shared split operator group (122) : array_obj_ref_1079_index_offset 
    ApIntAdd_group_122: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x0x_xlcssa_1078_scaled;
      array_obj_ref_1079_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1079_index_offset_req_0;
      array_obj_ref_1079_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1079_index_offset_req_1;
      array_obj_ref_1079_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_122_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_122_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_122",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 122
    -- shared split operator group (123) : array_obj_ref_1232_index_offset 
    ApIntAdd_group_123: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar412_1231_scaled;
      array_obj_ref_1232_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1232_index_offset_req_0;
      array_obj_ref_1232_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1232_index_offset_req_1;
      array_obj_ref_1232_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_123_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_123_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_123",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 123
    -- shared split operator group (124) : array_obj_ref_1552_index_offset 
    ApIntAdd_group_124: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1551_scaled;
      array_obj_ref_1552_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1552_index_offset_req_0;
      array_obj_ref_1552_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1552_index_offset_req_1;
      array_obj_ref_1552_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_124_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_124_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_124",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 124
    -- shared split operator group (125) : array_obj_ref_763_index_offset 
    ApIntAdd_group_125: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar426_762_scaled;
      array_obj_ref_763_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_763_index_offset_req_0;
      array_obj_ref_763_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_763_index_offset_req_1;
      array_obj_ref_763_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_125_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_125_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_125",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 125
    -- unary operator type_cast_1196_inst
    process(tmp19_1193) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp19_1193, tmp_var);
      type_cast_1196_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1690_inst
    process(call229_1563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call229_1563, tmp_var);
      type_cast_1690_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1698_inst
    process(call284_1695) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call284_1695, tmp_var);
      type_cast_1698_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_664_inst
    process(mul82_660) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", mul82_660, tmp_var);
      type_cast_664_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_692_inst
    process(tmp418_689) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp418_689, tmp_var);
      type_cast_692_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_727_inst
    process(tmp27_724) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", tmp27_724, tmp_var);
      type_cast_727_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_900_store_0 ptr_deref_1083_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_900_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1083_store_0_req_0;
      ptr_deref_900_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1083_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_900_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1083_store_0_req_1;
      ptr_deref_900_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1083_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_900_word_address_0 & ptr_deref_1083_word_address_0;
      data_in <= ptr_deref_900_data_0 & ptr_deref_1083_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1556_store_0 ptr_deref_1369_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1556_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1369_store_0_req_0;
      ptr_deref_1556_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1369_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1556_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1369_store_0_req_1;
      ptr_deref_1556_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1369_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1556_word_address_0 & ptr_deref_1369_word_address_0;
      data_in <= ptr_deref_1556_data_0 & ptr_deref_1369_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_maxpool_input_pipe_507_inst RPIPE_maxpool_input_pipe_569_inst RPIPE_maxpool_input_pipe_519_inst RPIPE_maxpool_input_pipe_544_inst RPIPE_maxpool_input_pipe_582_inst RPIPE_maxpool_input_pipe_632_inst RPIPE_maxpool_input_pipe_607_inst RPIPE_maxpool_input_pipe_557_inst RPIPE_maxpool_input_pipe_532_inst RPIPE_maxpool_input_pipe_619_inst RPIPE_maxpool_input_pipe_594_inst RPIPE_maxpool_input_pipe_1487_inst RPIPE_maxpool_input_pipe_1236_inst RPIPE_maxpool_input_pipe_1249_inst RPIPE_maxpool_input_pipe_1267_inst RPIPE_maxpool_input_pipe_1285_inst RPIPE_maxpool_input_pipe_1303_inst RPIPE_maxpool_input_pipe_1321_inst RPIPE_maxpool_input_pipe_1339_inst RPIPE_maxpool_input_pipe_1357_inst RPIPE_maxpool_input_pipe_444_inst RPIPE_maxpool_input_pipe_457_inst RPIPE_maxpool_input_pipe_469_inst RPIPE_maxpool_input_pipe_482_inst RPIPE_maxpool_input_pipe_494_inst RPIPE_maxpool_input_pipe_767_inst RPIPE_maxpool_input_pipe_780_inst RPIPE_maxpool_input_pipe_798_inst RPIPE_maxpool_input_pipe_816_inst RPIPE_maxpool_input_pipe_834_inst RPIPE_maxpool_input_pipe_852_inst RPIPE_maxpool_input_pipe_870_inst RPIPE_maxpool_input_pipe_888_inst RPIPE_maxpool_input_pipe_1014_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(271 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 33 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 33 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 33 downto 0);
      signal guard_vector : std_logic_vector( 33 downto 0);
      constant outBUFs : IntegerArray(33 downto 0) := (33 => 1, 32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(33 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false, 33 => false);
      constant guardBuffering: IntegerArray(33 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2, 33 => 2);
      -- 
    begin -- 
      reqL_unguarded(33) <= RPIPE_maxpool_input_pipe_507_inst_req_0;
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_569_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_519_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_544_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_582_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_632_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_607_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_557_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_532_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_619_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_594_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_1487_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_1236_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_1249_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1267_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_1285_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1303_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1321_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1339_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1357_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_444_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_457_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_469_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_482_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_494_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_767_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_780_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_798_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_816_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_834_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_852_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_870_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_888_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1014_inst_req_0;
      RPIPE_maxpool_input_pipe_507_inst_ack_0 <= ackL_unguarded(33);
      RPIPE_maxpool_input_pipe_569_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_519_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_544_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_582_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_632_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_607_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_557_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_532_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_619_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_594_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_1487_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_1236_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_1249_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1267_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_1285_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1303_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1321_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1339_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1357_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_444_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_457_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_469_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_482_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_494_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_767_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_780_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_798_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_816_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_834_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_852_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_870_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_888_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1014_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(33) <= RPIPE_maxpool_input_pipe_507_inst_req_1;
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_569_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_519_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_544_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_582_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_632_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_607_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_557_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_532_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_619_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_594_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_1487_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_1236_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_1249_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1267_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_1285_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1303_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1321_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1339_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1357_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_444_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_457_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_469_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_482_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_494_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_767_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_780_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_798_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_816_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_834_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_852_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_870_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_888_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1014_inst_req_1;
      RPIPE_maxpool_input_pipe_507_inst_ack_1 <= ackR_unguarded(33);
      RPIPE_maxpool_input_pipe_569_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_519_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_544_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_582_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_632_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_607_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_557_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_532_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_619_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_594_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_1487_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_1236_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_1249_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1267_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_1285_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1303_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1321_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1339_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1357_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_444_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_457_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_469_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_482_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_494_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_767_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_780_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_798_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_816_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_834_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_852_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_870_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_888_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1014_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      guard_vector(33)  <=  '1';
      call21_508 <= data_out(271 downto 264);
      call46_570 <= data_out(263 downto 256);
      call26_520 <= data_out(255 downto 248);
      call36_545 <= data_out(247 downto 240);
      call51_583 <= data_out(239 downto 232);
      call71_633 <= data_out(231 downto 224);
      call61_608 <= data_out(223 downto 216);
      call41_558 <= data_out(215 downto 208);
      call31_533 <= data_out(207 downto 200);
      call66_620 <= data_out(199 downto 192);
      call56_595 <= data_out(191 downto 184);
      callx_xi359_1488 <= data_out(183 downto 176);
      call164_1237 <= data_out(175 downto 168);
      call168_1250 <= data_out(167 downto 160);
      call174_1268 <= data_out(159 downto 152);
      call180_1286 <= data_out(151 downto 144);
      call186_1304 <= data_out(143 downto 136);
      call192_1322 <= data_out(135 downto 128);
      call198_1340 <= data_out(127 downto 120);
      call204_1358 <= data_out(119 downto 112);
      call_445 <= data_out(111 downto 104);
      call2_458 <= data_out(103 downto 96);
      call6_470 <= data_out(95 downto 88);
      call11_483 <= data_out(87 downto 80);
      call16_495 <= data_out(79 downto 72);
      call89_768 <= data_out(71 downto 64);
      call93_781 <= data_out(63 downto 56);
      call99_799 <= data_out(55 downto 48);
      call105_817 <= data_out(47 downto 40);
      call111_835 <= data_out(39 downto 32);
      call117_853 <= data_out(31 downto 24);
      call123_871 <= data_out(23 downto 16);
      call129_889 <= data_out(15 downto 8);
      callx_xi_1015 <= data_out(7 downto 0);
      maxpool_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_0_gI", nreqs => 34, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_0", data_width => 8,  num_reqs => 34,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1798_inst WPIPE_maxpool_output_pipe_1780_inst WPIPE_maxpool_output_pipe_1786_inst WPIPE_maxpool_output_pipe_1783_inst WPIPE_maxpool_output_pipe_1801_inst WPIPE_maxpool_output_pipe_1789_inst WPIPE_maxpool_output_pipe_1578_inst WPIPE_maxpool_output_pipe_1582_inst WPIPE_maxpool_output_pipe_1792_inst WPIPE_maxpool_output_pipe_1795_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(79 downto 0);
      signal sample_req, sample_ack : BooleanArray( 9 downto 0);
      signal update_req, update_ack : BooleanArray( 9 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 9 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 9 downto 0);
      signal guard_vector : std_logic_vector( 9 downto 0);
      constant inBUFs : IntegerArray(9 downto 0) := (9 => 0, 8 => 0, 7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(9 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false);
      constant guardBuffering: IntegerArray(9 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2);
      -- 
    begin -- 
      sample_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1798_inst_req_0;
      sample_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1780_inst_req_0;
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1786_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1783_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1801_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1789_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1578_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1582_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1792_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1795_inst_req_0;
      WPIPE_maxpool_output_pipe_1798_inst_ack_0 <= sample_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1780_inst_ack_0 <= sample_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1786_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1783_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1801_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1789_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1578_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1582_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1792_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1795_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(9) <= WPIPE_maxpool_output_pipe_1798_inst_req_1;
      update_req_unguarded(8) <= WPIPE_maxpool_output_pipe_1780_inst_req_1;
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1786_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1783_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1801_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1789_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1578_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1582_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1792_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1795_inst_req_1;
      WPIPE_maxpool_output_pipe_1798_inst_ack_1 <= update_ack_unguarded(9);
      WPIPE_maxpool_output_pipe_1780_inst_ack_1 <= update_ack_unguarded(8);
      WPIPE_maxpool_output_pipe_1786_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1783_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1801_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1789_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1578_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1582_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1792_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1795_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      data_in <= conv299_1719 & conv335_1779 & conv323_1759 & conv329_1769 & conv293_1709 & conv317_1749 & type_cast_1580_wire_constant & type_cast_1584_wire_constant & conv311_1739 & conv305_1729;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 10, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 10, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_1575_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1575_inst_req_0;
      WPIPE_num_out_pipe_1575_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1575_inst_req_1;
      WPIPE_num_out_pipe_1575_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= mul249_1574;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1695_call call_stmt_1563_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1695_call_req_0;
      reqL_unguarded(0) <= call_stmt_1563_call_req_0;
      call_stmt_1695_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1563_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1695_call_req_1;
      reqR_unguarded(0) <= call_stmt_1563_call_req_1;
      call_stmt_1695_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1563_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call284_1695 <= data_out(127 downto 64);
      call229_1563 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1662_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1662_call_req_0;
      call_stmt_1662_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1662_call_req_1;
      call_stmt_1662_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= conv255_1655 & conv261_1659;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 128,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(127 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1669_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1669_call_req_0;
      call_stmt_1669_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1669_call_req_1;
      call_stmt_1669_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul236_1569 & add33_542 & sub_1591 & sub269_1597 & add23_517 & add13_492;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 96,
        owidth => 96,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(95 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4033_start: Boolean;
  signal convolve_CP_4033_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal n_out_count_1912_1840_buf_req_0 : boolean;
  signal W_next_sum_1911_delayed_1_0_1938_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1898_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1843_inst_ack_0 : boolean;
  signal slice_1924_inst_req_1 : boolean;
  signal slice_1928_inst_ack_0 : boolean;
  signal n_out_count_1912_1840_buf_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1850_inst_ack_1 : boolean;
  signal RPIPE_input_pipe1_1843_inst_req_1 : boolean;
  signal W_next_sum_1911_delayed_1_0_1938_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_1898_inst_req_0 : boolean;
  signal slice_1928_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1843_inst_ack_1 : boolean;
  signal slice_1928_inst_req_0 : boolean;
  signal slice_1924_inst_ack_1 : boolean;
  signal W_next_sum_1911_delayed_1_0_1938_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_1850_inst_req_1 : boolean;
  signal do_while_stmt_1826_branch_req_0 : boolean;
  signal slice_1928_inst_ack_1 : boolean;
  signal type_cast_1936_inst_req_0 : boolean;
  signal type_cast_1944_inst_req_0 : boolean;
  signal type_cast_1936_inst_ack_0 : boolean;
  signal type_cast_1944_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1898_inst_req_1 : boolean;
  signal type_cast_1944_inst_req_1 : boolean;
  signal SUB_u32_u32_1864_inst_req_0 : boolean;
  signal type_cast_1936_inst_req_1 : boolean;
  signal type_cast_1936_inst_ack_1 : boolean;
  signal type_cast_1944_inst_ack_1 : boolean;
  signal SUB_u32_u32_1864_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_1898_inst_ack_1 : boolean;
  signal n_out_count_1912_1840_buf_req_1 : boolean;
  signal n_out_count_1912_1840_buf_ack_1 : boolean;
  signal W_next_sum_1906_delayed_1_0_1930_inst_req_0 : boolean;
  signal W_next_sum_1906_delayed_1_0_1930_inst_ack_0 : boolean;
  signal SUB_u32_u32_1864_inst_req_1 : boolean;
  signal W_next_sum_1906_delayed_1_0_1930_inst_req_1 : boolean;
  signal do_while_stmt_1826_branch_ack_1 : boolean;
  signal do_while_stmt_1826_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1942_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1942_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1942_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1942_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1812_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1812_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1812_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1812_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1815_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1815_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1815_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1815_inst_ack_1 : boolean;
  signal phi_stmt_1828_req_1 : boolean;
  signal phi_stmt_1828_req_0 : boolean;
  signal phi_stmt_1828_ack_0 : boolean;
  signal nmycount_1891_1831_buf_req_0 : boolean;
  signal nmycount_1891_1831_buf_ack_0 : boolean;
  signal nmycount_1891_1831_buf_req_1 : boolean;
  signal nmycount_1891_1831_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_1843_inst_req_0 : boolean;
  signal slice_1924_inst_ack_0 : boolean;
  signal slice_1924_inst_req_0 : boolean;
  signal W_next_sum_1911_delayed_1_0_1938_inst_ack_1 : boolean;
  signal phi_stmt_1832_req_1 : boolean;
  signal phi_stmt_1832_req_0 : boolean;
  signal phi_stmt_1832_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1934_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1934_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1934_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1934_inst_req_0 : boolean;
  signal nacc_1883_1835_buf_req_0 : boolean;
  signal nacc_1883_1835_buf_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1850_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_1850_inst_req_0 : boolean;
  signal nacc_1883_1835_buf_req_1 : boolean;
  signal nacc_1883_1835_buf_ack_1 : boolean;
  signal W_next_sum_1906_delayed_1_0_1930_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1919_inst_ack_1 : boolean;
  signal WPIPE_input_done_pipe_1919_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_1919_inst_ack_0 : boolean;
  signal SUB_u32_u32_1864_inst_ack_1 : boolean;
  signal phi_stmt_1836_req_1 : boolean;
  signal WPIPE_input_done_pipe_1919_inst_req_0 : boolean;
  signal phi_stmt_1836_req_0 : boolean;
  signal phi_stmt_1836_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4033_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4033_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4033_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4033_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4033: Block -- control-path 
    signal convolve_CP_4033_elements: BooleanArray(127 downto 0);
    -- 
  begin -- 
    convolve_CP_4033_elements(0) <= convolve_CP_4033_start;
    convolve_CP_4033_symbol <= convolve_CP_4033_elements(1);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1810/$entry
      -- CP-element group 0: 	 branch_block_stmt_1810/branch_block_stmt_1810__entry__
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825__entry__
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/$entry
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Sample/rr
      -- 
    rr_4055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(0), ack => RPIPE_num_out_pipe_1812_inst_req_0); -- 
    rr_4069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(0), ack => RPIPE_size_pipe_1815_inst_req_0); -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	127 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1810/$exit
      -- CP-element group 1: 	 branch_block_stmt_1810/branch_block_stmt_1810__exit__
      -- CP-element group 1: 	 branch_block_stmt_1810/do_while_stmt_1826__exit__
      -- 
    convolve_CP_4033_elements(1) <= convolve_CP_4033_elements(127);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Update/cr
      -- 
    ra_4056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1812_inst_ack_0, ack => convolve_CP_4033_elements(2)); -- 
    cr_4060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(2), ack => RPIPE_num_out_pipe_1812_inst_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_num_out_pipe_1812_Update/ca
      -- 
    ca_4061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1812_inst_ack_1, ack => convolve_CP_4033_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_update_start_
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Update/cr
      -- 
    ra_4070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1815_inst_ack_0, ack => convolve_CP_4033_elements(4)); -- 
    cr_4074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(4), ack => RPIPE_size_pipe_1815_inst_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/RPIPE_size_pipe_1815_Update/ca
      -- 
    ca_4075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1815_inst_ack_1, ack => convolve_CP_4033_elements(5)); -- 
    -- CP-element group 6:  join  transition  place  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825__exit__
      -- CP-element group 6: 	 branch_block_stmt_1810/do_while_stmt_1826__entry__
      -- CP-element group 6: 	 branch_block_stmt_1810/assign_stmt_1813_to_assign_stmt_1825/$exit
      -- 
    convolve_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 27) := "convolve_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(3) & convolve_CP_4033_elements(5);
      gj_convolve_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826__entry__
      -- CP-element group 7: 	 branch_block_stmt_1810/do_while_stmt_1826/$entry
      -- 
    convolve_CP_4033_elements(7) <= convolve_CP_4033_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	127 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826__exit__
      -- 
    -- Element group convolve_CP_4033_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_back
      -- 
    -- Element group convolve_CP_4033_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	125 
    -- CP-element group 10: 	126 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1810/do_while_stmt_1826/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_exit/$entry
      -- 
    convolve_CP_4033_elements(10) <= convolve_CP_4033_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	124 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_body_done
      -- 
    convolve_CP_4033_elements(11) <= convolve_CP_4033_elements(124);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	24 
    -- CP-element group 12: 	43 
    -- CP-element group 12: 	62 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4033_elements(12) <= convolve_CP_4033_elements(9);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	45 
    -- CP-element group 13: 	64 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4033_elements(13) <= convolve_CP_4033_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	21 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	75 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	83 
    -- CP-element group 14: 	123 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_4033_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	123 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/condition_evaluated
      -- 
    condition_evaluated_4090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(15), ack => do_while_stmt_1826_branch_req_0); -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(19) & convolve_CP_4033_elements(123);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	37 
    -- CP-element group 16: 	56 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_sample_start__ps
      -- CP-element group 16: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(20) & convolve_CP_4033_elements(37) & convolve_CP_4033_elements(56) & convolve_CP_4033_elements(19);
      gj_convolve_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	22 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	76 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	84 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	37 
    -- CP-element group 17: 	56 
    -- CP-element group 17:  members (4) 
      -- CP-element group 17: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_sample_completed_
      -- 
    convolve_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(22) & convolve_CP_4033_elements(40) & convolve_CP_4033_elements(59);
      gj_convolve_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: 	38 
    -- CP-element group 18: 	57 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	60 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_update_start__ps
      -- 
    convolve_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(21) & convolve_CP_4033_elements(38) & convolve_CP_4033_elements(57);
      gj_convolve_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	23 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	61 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(23) & convolve_CP_4033_elements(42) & convolve_CP_4033_elements(61);
      gj_convolve_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: 	86 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_sample_start_
      -- 
    convolve_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(17) & convolve_CP_4033_elements(86);
      gj_convolve_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	14 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	103 
    -- CP-element group 21: 	114 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_update_start_
      -- 
    convolve_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(91) & convolve_CP_4033_elements(103) & convolve_CP_4033_elements(114);
      gj_convolve_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	17 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_sample_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	90 
    -- CP-element group 23: 	101 
    -- CP-element group 23: 	112 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_update_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	12 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_loopback_trigger
      -- 
    convolve_CP_4033_elements(24) <= convolve_CP_4033_elements(12);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_loopback_sample_req
      -- CP-element group 25: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_loopback_sample_req_ps
      -- 
    phi_stmt_1828_loopback_sample_req_4105_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1828_loopback_sample_req_4105_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(25), ack => phi_stmt_1828_req_1); -- 
    -- Element group convolve_CP_4033_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	13 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_entry_trigger
      -- 
    convolve_CP_4033_elements(26) <= convolve_CP_4033_elements(13);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_entry_sample_req
      -- CP-element group 27: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_entry_sample_req_ps
      -- 
    phi_stmt_1828_entry_sample_req_4108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1828_entry_sample_req_4108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(27), ack => phi_stmt_1828_req_0); -- 
    -- Element group convolve_CP_4033_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_phi_mux_ack
      -- CP-element group 28: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1828_phi_mux_ack_ps
      -- 
    phi_stmt_1828_phi_mux_ack_4111_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1828_ack_0, ack => convolve_CP_4033_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_sample_start__ps
      -- CP-element group 29: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_sample_completed_
      -- 
    -- Element group convolve_CP_4033_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_update_start__ps
      -- CP-element group 30: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_update_start_
      -- 
    -- Element group convolve_CP_4033_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_update_completed__ps
      -- 
    convolve_CP_4033_elements(31) <= convolve_CP_4033_elements(32);
    -- CP-element group 32:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	31 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_mcount_var_1830_update_completed_
      -- 
    -- Element group convolve_CP_4033_elements(32) is a control-delay.
    cp_element_32_delay: control_delay_element  generic map(name => " 32_delay", delay_value => 1)  port map(req => convolve_CP_4033_elements(30), ack => convolve_CP_4033_elements(32), clk => clk, reset =>reset);
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Sample/req
      -- 
    req_4132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(33), ack => nmycount_1891_1831_buf_req_0); -- 
    -- Element group convolve_CP_4033_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Update/req
      -- 
    req_4137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(34), ack => nmycount_1891_1831_buf_req_1); -- 
    -- Element group convolve_CP_4033_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Sample/ack
      -- 
    ack_4133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1891_1831_buf_ack_0, ack => convolve_CP_4033_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nmycount_1831_Update/ack
      -- 
    ack_4138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_1891_1831_buf_ack_1, ack => convolve_CP_4033_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	17 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	82 
    -- CP-element group 37: 	86 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	16 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_sample_start_
      -- 
    convolve_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(17) & convolve_CP_4033_elements(78) & convolve_CP_4033_elements(82) & convolve_CP_4033_elements(86);
      gj_convolve_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	95 
    -- CP-element group 38: 	99 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	18 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_update_start_
      -- 
    convolve_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(95) & convolve_CP_4033_elements(99);
      gj_convolve_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_sample_start__ps
      -- 
    convolve_CP_4033_elements(39) <= convolve_CP_4033_elements(16);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_sample_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_update_start__ps
      -- 
    convolve_CP_4033_elements(41) <= convolve_CP_4033_elements(18);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	19 
    -- CP-element group 42: 	93 
    -- CP-element group 42: 	97 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_update_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	12 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_loopback_trigger
      -- 
    convolve_CP_4033_elements(43) <= convolve_CP_4033_elements(12);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_loopback_sample_req_ps
      -- 
    phi_stmt_1832_loopback_sample_req_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1832_loopback_sample_req_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(44), ack => phi_stmt_1832_req_1); -- 
    -- Element group convolve_CP_4033_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	13 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_entry_trigger
      -- 
    convolve_CP_4033_elements(45) <= convolve_CP_4033_elements(13);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_entry_sample_req_ps
      -- 
    phi_stmt_1832_entry_sample_req_4152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1832_entry_sample_req_4152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(46), ack => phi_stmt_1832_req_0); -- 
    -- Element group convolve_CP_4033_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1832_phi_mux_ack_ps
      -- 
    phi_stmt_1832_phi_mux_ack_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1832_ack_0, ack => convolve_CP_4033_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_sample_completed_
      -- 
    -- Element group convolve_CP_4033_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_update_start_
      -- 
    -- Element group convolve_CP_4033_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_update_completed__ps
      -- 
    convolve_CP_4033_elements(50) <= convolve_CP_4033_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_acc_var_1834_update_completed_
      -- 
    -- Element group convolve_CP_4033_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => convolve_CP_4033_elements(49), ack => convolve_CP_4033_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Sample/req
      -- 
    req_4176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(52), ack => nacc_1883_1835_buf_req_0); -- 
    -- Element group convolve_CP_4033_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_update_start_
      -- CP-element group 53: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Update/req
      -- 
    req_4181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(53), ack => nacc_1883_1835_buf_req_1); -- 
    -- Element group convolve_CP_4033_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Sample/ack
      -- 
    ack_4177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1883_1835_buf_ack_0, ack => convolve_CP_4033_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_nacc_1835_Update/ack
      -- 
    ack_4182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc_1883_1835_buf_ack_1, ack => convolve_CP_4033_elements(55)); -- 
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	14 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	17 
    -- CP-element group 56: 	86 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	16 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_sample_start_
      -- 
    convolve_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(17) & convolve_CP_4033_elements(86);
      gj_convolve_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	88 
    -- CP-element group 57: 	91 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	18 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_update_start_
      -- 
    convolve_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(88) & convolve_CP_4033_elements(91);
      gj_convolve_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_sample_start__ps
      -- 
    convolve_CP_4033_elements(58) <= convolve_CP_4033_elements(16);
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_sample_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	18 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_update_start__ps
      -- 
    convolve_CP_4033_elements(60) <= convolve_CP_4033_elements(18);
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	19 
    -- CP-element group 61: 	87 
    -- CP-element group 61: 	90 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_update_completed__ps
      -- 
    -- Element group convolve_CP_4033_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	12 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_loopback_trigger
      -- 
    convolve_CP_4033_elements(62) <= convolve_CP_4033_elements(12);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_loopback_sample_req
      -- CP-element group 63: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_loopback_sample_req_ps
      -- 
    phi_stmt_1836_loopback_sample_req_4193_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1836_loopback_sample_req_4193_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(63), ack => phi_stmt_1836_req_1); -- 
    -- Element group convolve_CP_4033_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	13 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_entry_trigger
      -- 
    convolve_CP_4033_elements(64) <= convolve_CP_4033_elements(13);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_entry_sample_req
      -- CP-element group 65: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_entry_sample_req_ps
      -- 
    phi_stmt_1836_entry_sample_req_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1836_entry_sample_req_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(65), ack => phi_stmt_1836_req_0); -- 
    -- Element group convolve_CP_4033_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_phi_mux_ack
      -- CP-element group 66: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/phi_stmt_1836_phi_mux_ack_ps
      -- 
    phi_stmt_1836_phi_mux_ack_4199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1836_ack_0, ack => convolve_CP_4033_elements(66)); -- 
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_sample_start__ps
      -- CP-element group 67: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_sample_completed_
      -- 
    -- Element group convolve_CP_4033_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_update_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_update_start_
      -- 
    -- Element group convolve_CP_4033_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	70 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_update_completed__ps
      -- 
    convolve_CP_4033_elements(69) <= convolve_CP_4033_elements(70);
    -- CP-element group 70:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	69 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1839_update_completed_
      -- 
    -- Element group convolve_CP_4033_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convolve_CP_4033_elements(68), ack => convolve_CP_4033_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_sample_start__ps
      -- 
    req_4220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(71), ack => n_out_count_1912_1840_buf_req_0); -- 
    -- Element group convolve_CP_4033_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_update_start_
      -- CP-element group 72: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Update/req
      -- CP-element group 72: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_update_start__ps
      -- 
    req_4225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(72), ack => n_out_count_1912_1840_buf_req_1); -- 
    -- Element group convolve_CP_4033_elements(72) is bound as output of CP function.
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_sample_completed__ps
      -- 
    ack_4221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1912_1840_buf_ack_0, ack => convolve_CP_4033_elements(73)); -- 
    -- CP-element group 74:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_update_completed__ps
      -- CP-element group 74: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/R_n_out_count_1840_Update/ack
      -- 
    ack_4226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_out_count_1912_1840_buf_ack_1, ack => convolve_CP_4033_elements(74)); -- 
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	14 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	78 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_sample_start_
      -- CP-element group 75: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Sample/rr
      -- CP-element group 75: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Sample/$entry
      -- 
    rr_4235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(75), ack => RPIPE_input_pipe1_1843_inst_req_0); -- 
    convolve_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(78);
      gj_convolve_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	17 
    -- CP-element group 76: 	77 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	95 
    -- CP-element group 76: 	99 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Update/cr
      -- CP-element group 76: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_update_start_
      -- 
    cr_4240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(76), ack => RPIPE_input_pipe1_1843_inst_req_1); -- 
    convolve_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(17) & convolve_CP_4033_elements(77) & convolve_CP_4033_elements(95) & convolve_CP_4033_elements(99);
      gj_convolve_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	76 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Sample/ra
      -- CP-element group 77: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_sample_completed_
      -- CP-element group 77: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Sample/$exit
      -- 
    ra_4236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1843_inst_ack_0, ack => convolve_CP_4033_elements(77)); -- 
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	93 
    -- CP-element group 78: 	97 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: 	75 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Update/ca
      -- CP-element group 78: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_Update/$exit
      -- CP-element group 78: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_input_pipe1_1843_update_completed_
      -- 
    ca_4241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1843_inst_ack_1, ack => convolve_CP_4033_elements(78)); -- 
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	82 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_sample_start_
      -- CP-element group 79: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Sample/$entry
      -- CP-element group 79: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Sample/rr
      -- 
    rr_4249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(79), ack => RPIPE_kernel_pipe1_1850_inst_req_0); -- 
    convolve_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(82);
      gj_convolve_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: 	81 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	88 
    -- CP-element group 80: 	95 
    -- CP-element group 80: 	99 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Update/cr
      -- CP-element group 80: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_update_start_
      -- 
    cr_4254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(80), ack => RPIPE_kernel_pipe1_1850_inst_req_1); -- 
    convolve_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(17) & convolve_CP_4033_elements(81) & convolve_CP_4033_elements(88) & convolve_CP_4033_elements(95) & convolve_CP_4033_elements(99);
      gj_convolve_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Sample/ra
      -- 
    ra_4250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1850_inst_ack_0, ack => convolve_CP_4033_elements(81)); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	87 
    -- CP-element group 82: 	93 
    -- CP-element group 82: 	97 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	37 
    -- CP-element group 82: 	79 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Update/ca
      -- CP-element group 82: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/RPIPE_kernel_pipe1_1850_update_completed_
      -- 
    ca_4255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_1850_inst_ack_1, ack => convolve_CP_4033_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	14 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Sample/rr
      -- 
    rr_4263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(83), ack => SUB_u32_u32_1864_inst_req_0); -- 
    convolve_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(14) & convolve_CP_4033_elements(85);
      gj_convolve_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	17 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	91 
    -- CP-element group 84: 	103 
    -- CP-element group 84: 	114 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Update/cr
      -- 
    cr_4268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(84), ack => SUB_u32_u32_1864_inst_req_1); -- 
    convolve_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(17) & convolve_CP_4033_elements(91) & convolve_CP_4033_elements(103) & convolve_CP_4033_elements(114);
      gj_convolve_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Sample/ra
      -- 
    ra_4264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1864_inst_ack_0, ack => convolve_CP_4033_elements(85)); -- 
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	90 
    -- CP-element group 86: 	101 
    -- CP-element group 86: 	112 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	20 
    -- CP-element group 86: 	37 
    -- CP-element group 86: 	56 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/SUB_u32_u32_1864_Update/ca
      -- 
    ca_4269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_1864_inst_ack_1, ack => convolve_CP_4033_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	61 
    -- CP-element group 87: 	82 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	89 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_sample_start_
      -- 
    req_4277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(87), ack => WPIPE_kernel_pipe1_1898_inst_req_0); -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(61) & convolve_CP_4033_elements(82) & convolve_CP_4033_elements(89);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-successors 
    -- CP-element group 88: 	57 
    -- CP-element group 88: 	80 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Sample/ack
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Update/req
      -- 
    ack_4278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1898_inst_ack_0, ack => convolve_CP_4033_elements(88)); -- 
    req_4282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(88), ack => WPIPE_kernel_pipe1_1898_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	124 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	87 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_kernel_pipe1_1898_Update/ack
      -- 
    ack_4283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_1898_inst_ack_1, ack => convolve_CP_4033_elements(89)); -- 
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	23 
    -- CP-element group 90: 	61 
    -- CP-element group 90: 	86 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	92 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Sample/req
      -- 
    req_4291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(90), ack => WPIPE_input_done_pipe_1919_inst_req_0); -- 
    convolve_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(23) & convolve_CP_4033_elements(61) & convolve_CP_4033_elements(86) & convolve_CP_4033_elements(92);
      gj_convolve_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	57 
    -- CP-element group 91: 	84 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_sample_completed_
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_update_start_
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Update/req
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Sample/$exit
      -- 
    ack_4292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1919_inst_ack_0, ack => convolve_CP_4033_elements(91)); -- 
    req_4296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(91), ack => WPIPE_input_done_pipe_1919_inst_req_1); -- 
    -- CP-element group 92:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	124 
    -- CP-element group 92: marked-successors 
    -- CP-element group 92: 	90 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_update_completed_
      -- CP-element group 92: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Update/ack
      -- CP-element group 92: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_input_done_pipe_1919_Update/$exit
      -- 
    ack_4297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_1919_inst_ack_1, ack => convolve_CP_4033_elements(92)); -- 
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	42 
    -- CP-element group 93: 	78 
    -- CP-element group 93: 	82 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	95 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_sample_start_
      -- 
    rr_4305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(93), ack => slice_1924_inst_req_0); -- 
    convolve_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(42) & convolve_CP_4033_elements(78) & convolve_CP_4033_elements(82) & convolve_CP_4033_elements(95);
      gj_convolve_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	107 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_update_start_
      -- 
    cr_4310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(94), ack => slice_1924_inst_req_1); -- 
    convolve_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4033_elements(107);
      gj_convolve_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: marked-successors 
    -- CP-element group 95: 	38 
    -- CP-element group 95: 	76 
    -- CP-element group 95: 	80 
    -- CP-element group 95: 	93 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Sample/ra
      -- CP-element group 95: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_sample_completed_
      -- 
    ra_4306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1924_inst_ack_0, ack => convolve_CP_4033_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	105 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Update/ca
      -- CP-element group 96: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1924_update_completed_
      -- 
    ca_4311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1924_inst_ack_1, ack => convolve_CP_4033_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	42 
    -- CP-element group 97: 	78 
    -- CP-element group 97: 	82 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Sample/rr
      -- 
    rr_4319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(97), ack => slice_1928_inst_req_0); -- 
    convolve_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(42) & convolve_CP_4033_elements(78) & convolve_CP_4033_elements(82) & convolve_CP_4033_elements(99);
      gj_convolve_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	118 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_update_start_
      -- 
    cr_4324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(98), ack => slice_1928_inst_req_1); -- 
    convolve_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4033_elements(118);
      gj_convolve_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	38 
    -- CP-element group 99: 	76 
    -- CP-element group 99: 	80 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Sample/ra
      -- CP-element group 99: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_sample_completed_
      -- 
    ra_4320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1928_inst_ack_0, ack => convolve_CP_4033_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	116 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/slice_1928_Update/ca
      -- 
    ca_4325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_1928_inst_ack_1, ack => convolve_CP_4033_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	23 
    -- CP-element group 101: 	86 
    -- CP-element group 101: marked-predecessors 
    -- CP-element group 101: 	103 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Sample/req
      -- 
    req_4333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(101), ack => W_next_sum_1906_delayed_1_0_1930_inst_req_0); -- 
    convolve_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(23) & convolve_CP_4033_elements(86) & convolve_CP_4033_elements(103);
      gj_convolve_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	107 
    -- CP-element group 102: 	110 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Update/req
      -- 
    req_4338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(102), ack => W_next_sum_1906_delayed_1_0_1930_inst_req_1); -- 
    convolve_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(107) & convolve_CP_4033_elements(110);
      gj_convolve_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103: marked-successors 
    -- CP-element group 103: 	21 
    -- CP-element group 103: 	84 
    -- CP-element group 103: 	101 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Sample/ack
      -- 
    ack_4334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1906_delayed_1_0_1930_inst_ack_0, ack => convolve_CP_4033_elements(103)); -- 
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104: 	109 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1932_Update/ack
      -- 
    ack_4339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1906_delayed_1_0_1930_inst_ack_1, ack => convolve_CP_4033_elements(104)); -- 
    -- CP-element group 105:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	96 
    -- CP-element group 105: 	104 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	107 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_sample_start_
      -- 
    rr_4347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(105), ack => type_cast_1936_inst_req_0); -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(96) & convolve_CP_4033_elements(104) & convolve_CP_4033_elements(107);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	110 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_update_start_
      -- CP-element group 106: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Update/$entry
      -- CP-element group 106: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Update/cr
      -- 
    cr_4352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(106), ack => type_cast_1936_inst_req_1); -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4033_elements(110);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: marked-successors 
    -- CP-element group 107: 	94 
    -- CP-element group 107: 	102 
    -- CP-element group 107: 	105 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Sample/$exit
      -- CP-element group 107: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Sample/ra
      -- CP-element group 107: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_sample_completed_
      -- 
    ra_4348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1936_inst_ack_0, ack => convolve_CP_4033_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Update/$exit
      -- CP-element group 108: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1936_Update/ca
      -- 
    ca_4353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1936_inst_ack_1, ack => convolve_CP_4033_elements(108)); -- 
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	104 
    -- CP-element group 109: 	108 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	122 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Sample/req
      -- 
    req_4361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(109), ack => WPIPE_maxpool_output_pipe_1934_inst_req_0); -- 
    convolve_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(104) & convolve_CP_4033_elements(108) & convolve_CP_4033_elements(122);
      gj_convolve_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	102 
    -- CP-element group 110: 	106 
    -- CP-element group 110:  members (6) 
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_update_start_
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Update/req
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Update/$entry
      -- CP-element group 110: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Sample/ack
      -- 
    ack_4362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1934_inst_ack_0, ack => convolve_CP_4033_elements(110)); -- 
    req_4366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(110), ack => WPIPE_maxpool_output_pipe_1934_inst_req_1); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	120 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Update/ack
      -- CP-element group 111: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1934_Update/$exit
      -- 
    ack_4367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1934_inst_ack_1, ack => convolve_CP_4033_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	23 
    -- CP-element group 112: 	86 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	114 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_sample_start_
      -- 
    req_4375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(112), ack => W_next_sum_1911_delayed_1_0_1938_inst_req_0); -- 
    convolve_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(23) & convolve_CP_4033_elements(86) & convolve_CP_4033_elements(114);
      gj_convolve_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	118 
    -- CP-element group 113: 	121 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Update/req
      -- CP-element group 113: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_update_start_
      -- 
    req_4380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(113), ack => W_next_sum_1911_delayed_1_0_1938_inst_req_1); -- 
    convolve_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(118) & convolve_CP_4033_elements(121);
      gj_convolve_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	21 
    -- CP-element group 114: 	84 
    -- CP-element group 114: 	112 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_sample_completed_
      -- 
    ack_4376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1911_delayed_1_0_1938_inst_ack_0, ack => convolve_CP_4033_elements(114)); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	120 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_Update/ack
      -- CP-element group 115: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/assign_stmt_1940_update_completed_
      -- 
    ack_4381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_next_sum_1911_delayed_1_0_1938_inst_ack_1, ack => convolve_CP_4033_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	100 
    -- CP-element group 116: 	115 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Sample/rr
      -- 
    rr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(116), ack => type_cast_1944_inst_req_0); -- 
    convolve_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(100) & convolve_CP_4033_elements(115) & convolve_CP_4033_elements(118);
      gj_convolve_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	121 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_update_start_
      -- CP-element group 117: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Update/cr
      -- 
    cr_4394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(117), ack => type_cast_1944_inst_req_1); -- 
    convolve_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= convolve_CP_4033_elements(121);
      gj_convolve_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	98 
    -- CP-element group 118: 	113 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Sample/ra
      -- 
    ra_4390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_0, ack => convolve_CP_4033_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/type_cast_1944_Update/ca
      -- 
    ca_4395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1944_inst_ack_1, ack => convolve_CP_4033_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	111 
    -- CP-element group 120: 	115 
    -- CP-element group 120: 	119 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	121 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Sample/$entry
      -- CP-element group 120: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Sample/req
      -- 
    req_4403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(120), ack => WPIPE_maxpool_output_pipe_1942_inst_req_0); -- 
    convolve_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(111) & convolve_CP_4033_elements(115) & convolve_CP_4033_elements(119) & convolve_CP_4033_elements(122);
      gj_convolve_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	120 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	113 
    -- CP-element group 121: 	117 
    -- CP-element group 121:  members (6) 
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_update_start_
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Update/req
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Sample/ack
      -- CP-element group 121: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Sample/$exit
      -- 
    ack_4404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1942_inst_ack_0, ack => convolve_CP_4033_elements(121)); -- 
    req_4408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4033_elements(121), ack => WPIPE_maxpool_output_pipe_1942_inst_req_1); -- 
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	109 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Update/ack
      -- CP-element group 122: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/WPIPE_maxpool_output_pipe_1942_Update/$exit
      -- 
    ack_4409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1942_inst_ack_1, ack => convolve_CP_4033_elements(122)); -- 
    -- CP-element group 123:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	14 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	15 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4033_elements(123) is a control-delay.
    cp_element_123_delay: control_delay_element  generic map(name => " 123_delay", delay_value => 1)  port map(req => convolve_CP_4033_elements(14), ack => convolve_CP_4033_elements(123), clk => clk, reset =>reset);
    -- CP-element group 124:  join  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	89 
    -- CP-element group 124: 	92 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	11 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1810/do_while_stmt_1826/do_while_stmt_1826_loop_body/$exit
      -- 
    convolve_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4033_elements(89) & convolve_CP_4033_elements(92) & convolve_CP_4033_elements(122);
      gj_convolve_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4033_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	10 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (2) 
      -- CP-element group 125: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_exit/ack
      -- CP-element group 125: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_exit/$exit
      -- 
    ack_4414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1826_branch_ack_0, ack => convolve_CP_4033_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	10 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (2) 
      -- CP-element group 126: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_taken/ack
      -- CP-element group 126: 	 branch_block_stmt_1810/do_while_stmt_1826/loop_taken/$exit
      -- 
    ack_4418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1826_branch_ack_1, ack => convolve_CP_4033_elements(126)); -- 
    -- CP-element group 127:  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	8 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	1 
    -- CP-element group 127:  members (1) 
      -- CP-element group 127: 	 branch_block_stmt_1810/do_while_stmt_1826/$exit
      -- 
    convolve_CP_4033_elements(127) <= convolve_CP_4033_elements(8);
    convolve_do_while_stmt_1826_terminator_4419: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1826_terminator_4419", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4033_elements(11),loop_continue => convolve_CP_4033_elements(126),loop_terminate => convolve_CP_4033_elements(125),loop_back => convolve_CP_4033_elements(9),loop_exit => convolve_CP_4033_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1828_phi_seq_4139_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4033_elements(26);
      convolve_CP_4033_elements(29)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4033_elements(29);
      convolve_CP_4033_elements(30)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4033_elements(31);
      convolve_CP_4033_elements(27) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4033_elements(24);
      convolve_CP_4033_elements(33)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4033_elements(35);
      convolve_CP_4033_elements(34)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4033_elements(36);
      convolve_CP_4033_elements(25) <= phi_mux_reqs(1);
      phi_stmt_1828_phi_seq_4139 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1828_phi_seq_4139") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4033_elements(16), 
          phi_sample_ack => convolve_CP_4033_elements(22), 
          phi_update_req => convolve_CP_4033_elements(18), 
          phi_update_ack => convolve_CP_4033_elements(23), 
          phi_mux_ack => convolve_CP_4033_elements(28), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1832_phi_seq_4183_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4033_elements(45);
      convolve_CP_4033_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4033_elements(48);
      convolve_CP_4033_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4033_elements(50);
      convolve_CP_4033_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4033_elements(43);
      convolve_CP_4033_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4033_elements(54);
      convolve_CP_4033_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4033_elements(55);
      convolve_CP_4033_elements(44) <= phi_mux_reqs(1);
      phi_stmt_1832_phi_seq_4183 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1832_phi_seq_4183") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4033_elements(39), 
          phi_sample_ack => convolve_CP_4033_elements(40), 
          phi_update_req => convolve_CP_4033_elements(41), 
          phi_update_ack => convolve_CP_4033_elements(42), 
          phi_mux_ack => convolve_CP_4033_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1836_phi_seq_4227_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4033_elements(64);
      convolve_CP_4033_elements(67)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4033_elements(67);
      convolve_CP_4033_elements(68)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4033_elements(69);
      convolve_CP_4033_elements(65) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4033_elements(62);
      convolve_CP_4033_elements(71)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4033_elements(73);
      convolve_CP_4033_elements(72)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4033_elements(74);
      convolve_CP_4033_elements(63) <= phi_mux_reqs(1);
      phi_stmt_1836_phi_seq_4227 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1836_phi_seq_4227") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4033_elements(58), 
          phi_sample_ack => convolve_CP_4033_elements(59), 
          phi_update_req => convolve_CP_4033_elements(60), 
          phi_update_ack => convolve_CP_4033_elements(61), 
          phi_mux_ack => convolve_CP_4033_elements(66), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4091_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4033_elements(12);
        preds(1)  <= convolve_CP_4033_elements(13);
        entry_tmerge_4091 : transition_merge -- 
          generic map(name => " entry_tmerge_4091")
          port map (preds => preds, symbol_out => convolve_CP_4033_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_1908_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_1889_wire : std_logic_vector(31 downto 0);
    signal MUX_1909_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_1844_1844_delayed_1_0_1865 : std_logic_vector(31 downto 0);
    signal acc_1832 : std_logic_vector(15 downto 0);
    signal acc_val_1877 : std_logic_vector(15 downto 0);
    signal acc_val_dn_1929 : std_logic_vector(7 downto 0);
    signal acc_val_up_1925 : std_logic_vector(7 downto 0);
    signal acc_var_1825 : std_logic_vector(15 downto 0);
    signal all_done_flag_1917 : std_logic_vector(0 downto 0);
    signal iread_1844 : std_logic_vector(15 downto 0);
    signal ival_1848 : std_logic_vector(15 downto 0);
    signal konst_1863_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1880_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1886_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1888_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1920_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1947_wire_constant : std_logic_vector(0 downto 0);
    signal kread_1851 : std_logic_vector(15 downto 0);
    signal kval_1855 : std_logic_vector(15 downto 0);
    signal mcount_var_1820 : std_logic_vector(31 downto 0);
    signal mul_val_1860 : std_logic_vector(15 downto 0);
    signal mycount_1828 : std_logic_vector(31 downto 0);
    signal n_out_count_1912 : std_logic_vector(15 downto 0);
    signal n_out_count_1912_1840_buffered : std_logic_vector(15 downto 0);
    signal nacc_1883 : std_logic_vector(15 downto 0);
    signal nacc_1883_1835_buffered : std_logic_vector(15 downto 0);
    signal next_sum_1870 : std_logic_vector(0 downto 0);
    signal next_sum_1906_delayed_1_0_1932 : std_logic_vector(0 downto 0);
    signal next_sum_1911_delayed_1_0_1940 : std_logic_vector(0 downto 0);
    signal nmycount_1891 : std_logic_vector(31 downto 0);
    signal nmycount_1891_1831_buffered : std_logic_vector(31 downto 0);
    signal num_out_1813 : std_logic_vector(15 downto 0);
    signal out_count_1836 : std_logic_vector(15 downto 0);
    signal out_done_flag_1896 : std_logic_vector(0 downto 0);
    signal size_1816 : std_logic_vector(31 downto 0);
    signal type_cast_1839_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1873_wire : std_logic_vector(15 downto 0);
    signal type_cast_1875_wire : std_logic_vector(15 downto 0);
    signal type_cast_1905_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1936_wire : std_logic_vector(7 downto 0);
    signal type_cast_1944_wire : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    acc_var_1825 <= "0000000000000000";
    konst_1863_wire_constant <= "00000000000000000000000000000001";
    konst_1880_wire_constant <= "0000000000000000";
    konst_1886_wire_constant <= "00000000000000000000000000000000";
    konst_1888_wire_constant <= "00000000000000000000000000000001";
    konst_1907_wire_constant <= "0000000000000001";
    konst_1920_wire_constant <= "1";
    konst_1947_wire_constant <= "1";
    mcount_var_1820 <= "00000000000000000000000000000000";
    type_cast_1839_wire_constant <= "0000000000000001";
    type_cast_1905_wire_constant <= "0000000000000001";
    phi_stmt_1828: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= mcount_var_1820 & nmycount_1891_1831_buffered;
      req <= phi_stmt_1828_req_0 & phi_stmt_1828_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1828",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1828_ack_0,
          idata => idata,
          odata => mycount_1828,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1828
    phi_stmt_1832: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= acc_var_1825 & nacc_1883_1835_buffered;
      req <= phi_stmt_1832_req_0 & phi_stmt_1832_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1832",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1832_ack_0,
          idata => idata,
          odata => acc_1832,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1832
    phi_stmt_1836: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1839_wire_constant & n_out_count_1912_1840_buffered;
      req <= phi_stmt_1836_req_0 & phi_stmt_1836_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1836",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1836_ack_0,
          idata => idata,
          odata => out_count_1836,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1836
    -- flow-through select operator MUX_1882_inst
    nacc_1883 <= konst_1880_wire_constant when (next_sum_1870(0) /=  '0') else acc_val_1877;
    -- flow-through select operator MUX_1890_inst
    nmycount_1891 <= konst_1886_wire_constant when (next_sum_1870(0) /=  '0') else ADD_u32_u32_1889_wire;
    -- flow-through select operator MUX_1909_inst
    MUX_1909_wire <= type_cast_1905_wire_constant when (out_done_flag_1896(0) /=  '0') else ADD_u16_u16_1908_wire;
    -- flow-through select operator MUX_1911_inst
    n_out_count_1912 <= MUX_1909_wire when (next_sum_1870(0) /=  '0') else out_count_1836;
    slice_1924_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1924_inst_req_0;
      slice_1924_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1924_inst_req_1;
      slice_1924_inst_ack_1<= update_ack(0);
      slice_1924_inst: SliceSplitProtocol generic map(name => "slice_1924_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1877, dout => acc_val_up_1925, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_1928_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_1928_inst_req_0;
      slice_1928_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_1928_inst_req_1;
      slice_1928_inst_ack_1<= update_ack(0);
      slice_1928_inst: SliceSplitProtocol generic map(name => "slice_1928_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => acc_val_1877, dout => acc_val_dn_1929, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_next_sum_1906_delayed_1_0_1930_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1906_delayed_1_0_1930_inst_req_0;
      W_next_sum_1906_delayed_1_0_1930_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1906_delayed_1_0_1930_inst_req_1;
      W_next_sum_1906_delayed_1_0_1930_inst_ack_1<= rack(0);
      W_next_sum_1906_delayed_1_0_1930_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1906_delayed_1_0_1930_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1870,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1906_delayed_1_0_1932,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_next_sum_1911_delayed_1_0_1938_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_next_sum_1911_delayed_1_0_1938_inst_req_0;
      W_next_sum_1911_delayed_1_0_1938_inst_ack_0<= wack(0);
      rreq(0) <= W_next_sum_1911_delayed_1_0_1938_inst_req_1;
      W_next_sum_1911_delayed_1_0_1938_inst_ack_1<= rack(0);
      W_next_sum_1911_delayed_1_0_1938_inst : InterlockBuffer generic map ( -- 
        name => "W_next_sum_1911_delayed_1_0_1938_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => next_sum_1870,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => next_sum_1911_delayed_1_0_1940,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_out_count_1912_1840_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_out_count_1912_1840_buf_req_0;
      n_out_count_1912_1840_buf_ack_0<= wack(0);
      rreq(0) <= n_out_count_1912_1840_buf_req_1;
      n_out_count_1912_1840_buf_ack_1<= rack(0);
      n_out_count_1912_1840_buf : InterlockBuffer generic map ( -- 
        name => "n_out_count_1912_1840_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_out_count_1912,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_out_count_1912_1840_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc_1883_1835_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc_1883_1835_buf_req_0;
      nacc_1883_1835_buf_ack_0<= wack(0);
      rreq(0) <= nacc_1883_1835_buf_req_1;
      nacc_1883_1835_buf_ack_1<= rack(0);
      nacc_1883_1835_buf : InterlockBuffer generic map ( -- 
        name => "nacc_1883_1835_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc_1883,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc_1883_1835_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_1891_1831_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_1891_1831_buf_req_0;
      nmycount_1891_1831_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_1891_1831_buf_req_1;
      nmycount_1891_1831_buf_ack_1<= rack(0);
      nmycount_1891_1831_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_1891_1831_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_1891,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_1891_1831_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1847_inst
    process(iread_1844) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := iread_1844(15 downto 0);
      ival_1848 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1854_inst
    process(kread_1851) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := kread_1851(15 downto 0);
      kval_1855 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1873_inst
    process(acc_1832) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := acc_1832(15 downto 0);
      type_cast_1873_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1875_inst
    process(mul_val_1860) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := mul_val_1860(15 downto 0);
      type_cast_1875_wire <= tmp_var; -- 
    end process;
    type_cast_1936_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1936_inst_req_0;
      type_cast_1936_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1936_inst_req_1;
      type_cast_1936_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1906_delayed_1_0_1932(0);
      type_cast_1936_inst_gI: SplitGuardInterface generic map(name => "type_cast_1936_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1936_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1936_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_up_1925,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1936_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1944_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1944_inst_req_0;
      type_cast_1944_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1944_inst_req_1;
      type_cast_1944_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  next_sum_1911_delayed_1_0_1940(0);
      type_cast_1944_inst_gI: SplitGuardInterface generic map(name => "type_cast_1944_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1944_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1944_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc_val_dn_1929,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1944_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1826_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_1947_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1826_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1826_branch_req_0,
          ack0 => do_while_stmt_1826_branch_ack_0,
          ack1 => do_while_stmt_1826_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i16_i16_1876_inst
    process(type_cast_1873_wire, type_cast_1875_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_1873_wire, type_cast_1875_wire, tmp_var);
      acc_val_1877 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1908_inst
    process(out_count_1836) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(out_count_1836, konst_1907_wire_constant, tmp_var);
      ADD_u16_u16_1908_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1889_inst
    process(mycount_1828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_1828, konst_1888_wire_constant, tmp_var);
      ADD_u32_u32_1889_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1916_inst
    process(out_done_flag_1896, next_sum_1870) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_1896, next_sum_1870, tmp_var);
      all_done_flag_1917 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_1895_inst
    process(out_count_1836, num_out_1813) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(out_count_1836, num_out_1813, tmp_var);
      out_done_flag_1896 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1869_inst
    process(mycount_1828, SUB_u32_u32_1844_1844_delayed_1_0_1865) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycount_1828, SUB_u32_u32_1844_1844_delayed_1_0_1865, tmp_var);
      next_sum_1870 <= tmp_var; --
    end process;
    -- binary operator MUL_i16_i16_1859_inst
    process(kval_1855, ival_1848) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval_1855, ival_1848, tmp_var);
      mul_val_1860 <= tmp_var; --
    end process;
    -- shared split operator group (7) : SUB_u32_u32_1864_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= size_1816;
      SUB_u32_u32_1844_1844_delayed_1_0_1865 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_1864_inst_req_0;
      SUB_u32_u32_1864_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_1864_inst_req_1;
      SUB_u32_u32_1864_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared inport operator group (0) : RPIPE_input_pipe1_1843_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1843_inst_req_0;
      RPIPE_input_pipe1_1843_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1843_inst_req_1;
      RPIPE_input_pipe1_1843_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      iread_1844 <= data_out(15 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_kernel_pipe1_1850_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_1850_inst_req_0;
      RPIPE_kernel_pipe1_1850_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_1850_inst_req_1;
      RPIPE_kernel_pipe1_1850_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      kread_1851 <= data_out(15 downto 0);
      kernel_pipe1_read_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_1: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_num_out_pipe_1812_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1812_inst_req_0;
      RPIPE_num_out_pipe_1812_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1812_inst_req_1;
      RPIPE_num_out_pipe_1812_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      num_out_1813 <= data_out(15 downto 0);
      num_out_pipe_read_2_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_2: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_size_pipe_1815_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1815_inst_req_0;
      RPIPE_size_pipe_1815_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1815_inst_req_1;
      RPIPE_size_pipe_1815_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      size_1816 <= data_out(31 downto 0);
      size_pipe_read_3_gI: SplitGuardInterface generic map(name => "size_pipe_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_3: InputPortRevised -- 
        generic map ( name => "size_pipe_read_3", data_width => 32,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_input_done_pipe_1919_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_1919_inst_req_0;
      WPIPE_input_done_pipe_1919_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_1919_inst_req_1;
      WPIPE_input_done_pipe_1919_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= all_done_flag_1917(0);
      data_in <= konst_1920_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe1_1898_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_1898_inst_req_0;
      WPIPE_kernel_pipe1_1898_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_1898_inst_req_1;
      WPIPE_kernel_pipe1_1898_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  not out_done_flag_1896(0);
      data_in <= kread_1851;
      kernel_pipe1_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_maxpool_output_pipe_1934_inst WPIPE_maxpool_output_pipe_1942_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1934_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1942_inst_req_0;
      WPIPE_maxpool_output_pipe_1934_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1942_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1934_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1942_inst_req_1;
      WPIPE_maxpool_output_pipe_1934_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1942_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= next_sum_1911_delayed_1_0_1940(0);
      guard_vector(1)  <= next_sum_1906_delayed_1_0_1932(0);
      data_in <= type_cast_1936_wire & type_cast_1944_wire;
      maxpool_output_pipe_write_2_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 2, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(63 downto 0);
    end_add : in  std_logic_vector(63 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 128)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(63 downto 0);
  signal start_add_update_enable: Boolean;
  signal end_add_buffer :  std_logic_vector(63 downto 0);
  signal end_add_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_671_start: Boolean;
  signal loadKernelChannel_CP_671_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_437_inst_req_1 : boolean;
  signal type_cast_437_inst_ack_1 : boolean;
  signal phi_stmt_361_req_1 : boolean;
  signal my_fetch_344_364_buf_ack_0 : boolean;
  signal phi_stmt_361_req_0 : boolean;
  signal ptr_deref_411_load_0_req_1 : boolean;
  signal phi_stmt_361_ack_0 : boolean;
  signal WPIPE_size_pipe_433_inst_req_1 : boolean;
  signal addr_of_403_final_reg_req_0 : boolean;
  signal ptr_deref_411_load_0_ack_1 : boolean;
  signal addr_of_403_final_reg_ack_0 : boolean;
  signal type_cast_437_inst_req_0 : boolean;
  signal WPIPE_size_pipe_433_inst_ack_1 : boolean;
  signal nfetch_val_424_363_buf_ack_0 : boolean;
  signal my_fetch_344_364_buf_req_1 : boolean;
  signal my_fetch_344_364_buf_req_0 : boolean;
  signal addr_of_403_final_reg_req_1 : boolean;
  signal addr_of_403_final_reg_ack_1 : boolean;
  signal my_fetch_344_364_buf_ack_1 : boolean;
  signal W_fn_399_delayed_13_0_413_inst_ack_0 : boolean;
  signal do_while_stmt_355_branch_ack_0 : boolean;
  signal W_fetch_val_401_delayed_13_0_416_inst_req_1 : boolean;
  signal WPIPE_size_pipe_433_inst_ack_0 : boolean;
  signal type_cast_437_inst_ack_0 : boolean;
  signal W_fn_399_delayed_13_0_413_inst_req_1 : boolean;
  signal W_fn_399_delayed_13_0_413_inst_req_0 : boolean;
  signal WPIPE_size_pipe_433_inst_req_0 : boolean;
  signal W_fetch_val_401_delayed_13_0_416_inst_req_0 : boolean;
  signal nfetch_val_424_363_buf_req_0 : boolean;
  signal nfetch_val_424_363_buf_req_1 : boolean;
  signal W_fn_393_delayed_7_0_405_inst_req_0 : boolean;
  signal W_fn_393_delayed_7_0_405_inst_ack_0 : boolean;
  signal W_fn_399_delayed_13_0_413_inst_ack_1 : boolean;
  signal W_fetch_val_401_delayed_13_0_416_inst_ack_0 : boolean;
  signal nfetch_val_424_363_buf_ack_1 : boolean;
  signal do_while_stmt_355_branch_ack_1 : boolean;
  signal array_obj_ref_402_index_offset_req_0 : boolean;
  signal array_obj_ref_402_index_offset_ack_0 : boolean;
  signal array_obj_ref_402_index_offset_req_1 : boolean;
  signal W_fn_393_delayed_7_0_405_inst_req_1 : boolean;
  signal array_obj_ref_402_index_offset_ack_1 : boolean;
  signal W_fn_393_delayed_7_0_405_inst_ack_1 : boolean;
  signal ptr_deref_411_load_0_ack_0 : boolean;
  signal ptr_deref_411_load_0_req_0 : boolean;
  signal array_obj_ref_338_index_offset_req_0 : boolean;
  signal array_obj_ref_338_index_offset_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_386_inst_ack_1 : boolean;
  signal array_obj_ref_338_index_offset_req_1 : boolean;
  signal array_obj_ref_338_index_offset_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_386_inst_req_1 : boolean;
  signal addr_of_339_final_reg_req_0 : boolean;
  signal addr_of_339_final_reg_ack_0 : boolean;
  signal addr_of_339_final_reg_req_1 : boolean;
  signal addr_of_339_final_reg_ack_1 : boolean;
  signal WPIPE_kernel_pipe1_386_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_386_inst_req_0 : boolean;
  signal ptr_deref_343_load_0_req_0 : boolean;
  signal ptr_deref_343_load_0_ack_0 : boolean;
  signal start_add_360_buf_ack_1 : boolean;
  signal ptr_deref_343_load_0_req_1 : boolean;
  signal ptr_deref_343_load_0_ack_1 : boolean;
  signal W_fetch_val_401_delayed_13_0_416_inst_ack_1 : boolean;
  signal start_add_360_buf_req_1 : boolean;
  signal RPIPE_input_done_pipe_352_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_352_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_352_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_352_inst_ack_1 : boolean;
  signal do_while_stmt_355_branch_req_0 : boolean;
  signal phi_stmt_357_req_0 : boolean;
  signal phi_stmt_357_req_1 : boolean;
  signal phi_stmt_357_ack_0 : boolean;
  signal nmycount_379_359_buf_req_0 : boolean;
  signal nmycount_379_359_buf_ack_0 : boolean;
  signal nmycount_379_359_buf_req_1 : boolean;
  signal nmycount_379_359_buf_ack_1 : boolean;
  signal start_add_360_buf_req_0 : boolean;
  signal start_add_360_buf_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 128) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(63 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(63 downto 0);
  in_buffer_data_in(127 downto 64) <= end_add;
  end_add_buffer <= in_buffer_data_out(127 downto 64);
  in_buffer_data_in(tag_length + 127 downto 128) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 127 downto 128);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_671_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_671_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_671: Block -- control-path 
    signal loadKernelChannel_CP_671_elements: BooleanArray(94 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_671_elements(0) <= loadKernelChannel_CP_671_start;
    loadKernelChannel_CP_671_symbol <= loadKernelChannel_CP_671_elements(94);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	6 
    -- CP-element group 0:  members (29) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_update_start_
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_resized_1
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_scaled_1
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_computed_1
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_resize_1/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_resize_1/$exit
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_resize_1/index_resize_req
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_resize_1/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_scale_1/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_scale_1/$exit
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_scale_1/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_index_scale_1/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_update_start
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Sample/req
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Update/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Update/req
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_complete/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_complete/req
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_update_start_
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_sample_start_
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Sample/rr
      -- 
    req_721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => addr_of_339_final_reg_req_1); -- 
    req_701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_338_index_offset_req_0); -- 
    cr_766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => ptr_deref_343_load_0_req_1); -- 
    req_706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => array_obj_ref_338_index_offset_req_1); -- 
    rr_780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(0), ack => RPIPE_input_done_pipe_352_inst_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	9 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_sample_complete
      -- CP-element group 1: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Sample/ack
      -- 
    ack_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_338_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (11) 
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_sample_start_
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_root_address_calculated
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_offset_calculated
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Update/$exit
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_final_index_sum_regn_Update/ack
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_base_plus_offset/$entry
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_base_plus_offset/$exit
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/array_obj_ref_338_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_request/$entry
      -- CP-element group 2: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_request/req
      -- 
    ack_707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_338_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(2)); -- 
    req_716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(2), ack => addr_of_339_final_reg_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_sample_completed_
      -- CP-element group 3: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_request/$exit
      -- CP-element group 3: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_request/ack
      -- 
    ack_717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_339_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (24) 
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_update_completed_
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_complete/$exit
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/addr_of_339_complete/ack
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_sample_start_
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_address_calculated
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_word_address_calculated
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_root_address_calculated
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_address_resized
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_addr_resize/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_addr_resize/$exit
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_addr_resize/base_resize_req
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_addr_resize/base_resize_ack
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_plus_offset/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_plus_offset/$exit
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_plus_offset/sum_rename_req
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_base_plus_offset/sum_rename_ack
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_word_addrgen/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_word_addrgen/$exit
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_word_addrgen/root_register_req
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_word_addrgen/root_register_ack
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/word_0/$entry
      -- CP-element group 4: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/word_0/rr
      -- 
    ack_722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_339_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(4)); -- 
    rr_755_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_755_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(4), ack => ptr_deref_343_load_0_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_sample_completed_
      -- CP-element group 5: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/$exit
      -- CP-element group 5: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/$exit
      -- CP-element group 5: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Sample/word_access_start/word_0/ra
      -- 
    ra_756_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_update_completed_
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/$exit
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/$exit
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/ptr_deref_343_Merge/$entry
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/ptr_deref_343_Merge/$exit
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/ptr_deref_343_Merge/merge_req
      -- CP-element group 6: 	 assign_stmt_333_to_assign_stmt_353/ptr_deref_343_Update/ptr_deref_343_Merge/merge_ack
      -- 
    ca_767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_343_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_sample_completed_
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_update_start_
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Sample/ra
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Update/$entry
      -- CP-element group 7: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Update/cr
      -- 
    ra_781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_352_inst_ack_0, ack => loadKernelChannel_CP_671_elements(7)); -- 
    cr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(7), ack => RPIPE_input_done_pipe_352_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_update_completed_
      -- CP-element group 8: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Update/$exit
      -- CP-element group 8: 	 assign_stmt_333_to_assign_stmt_353/RPIPE_input_done_pipe_352_Update/ca
      -- 
    ca_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_352_inst_ack_1, ack => loadKernelChannel_CP_671_elements(8)); -- 
    -- CP-element group 9:  join  transition  place  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	1 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (4) 
      -- CP-element group 9: 	 assign_stmt_333_to_assign_stmt_353/$exit
      -- CP-element group 9: 	 branch_block_stmt_354/$entry
      -- CP-element group 9: 	 branch_block_stmt_354/branch_block_stmt_354__entry__
      -- CP-element group 9: 	 branch_block_stmt_354/do_while_stmt_355__entry__
      -- 
    loadKernelChannel_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "loadKernelChannel_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(1) & loadKernelChannel_CP_671_elements(8) & loadKernelChannel_CP_671_elements(6);
      gj_loadKernelChannel_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  place  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	90 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	91 
    -- CP-element group 10: 	92 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_Update/cr
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_438/$entry
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_Sample/rr
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_Update/$entry
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_sample_start_
      -- CP-element group 10: 	 assign_stmt_438/type_cast_437_update_start_
      -- CP-element group 10: 	 branch_block_stmt_354/$exit
      -- CP-element group 10: 	 branch_block_stmt_354/branch_block_stmt_354__exit__
      -- CP-element group 10: 	 branch_block_stmt_354/do_while_stmt_355__exit__
      -- 
    cr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => type_cast_437_inst_req_1); -- 
    rr_1094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(10), ack => type_cast_437_inst_req_0); -- 
    loadKernelChannel_CP_671_elements(10) <= loadKernelChannel_CP_671_elements(90);
    -- CP-element group 11:  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_354/do_while_stmt_355/$entry
      -- CP-element group 11: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355__entry__
      -- 
    loadKernelChannel_CP_671_elements(11) <= loadKernelChannel_CP_671_elements(9);
    -- CP-element group 12:  merge  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	90 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355__exit__
      -- 
    -- Element group loadKernelChannel_CP_671_elements(12) is bound as output of CP function.
    -- CP-element group 13:  merge  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	16 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_354/do_while_stmt_355/loop_back
      -- 
    -- Element group loadKernelChannel_CP_671_elements(13) is bound as output of CP function.
    -- CP-element group 14:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	88 
    -- CP-element group 14: 	89 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_354/do_while_stmt_355/loop_exit/$entry
      -- CP-element group 14: 	 branch_block_stmt_354/do_while_stmt_355/loop_taken/$entry
      -- CP-element group 14: 	 branch_block_stmt_354/do_while_stmt_355/condition_done
      -- 
    loadKernelChannel_CP_671_elements(14) <= loadKernelChannel_CP_671_elements(19);
    -- CP-element group 15:  branch  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	87 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_354/do_while_stmt_355/loop_body_done
      -- 
    loadKernelChannel_CP_671_elements(15) <= loadKernelChannel_CP_671_elements(87);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	13 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	28 
    -- CP-element group 16: 	47 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_671_elements(16) <= loadKernelChannel_CP_671_elements(13);
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	49 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_671_elements(17) <= loadKernelChannel_CP_671_elements(11);
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	86 
    -- CP-element group 18: 	25 
    -- CP-element group 18: 	41 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	64 
    -- CP-element group 18: 	65 
    -- CP-element group 18: 	24 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/$entry
      -- CP-element group 18: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(18) is bound as output of CP function.
    -- CP-element group 19:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	86 
    -- CP-element group 19: 	27 
    -- CP-element group 19: 	23 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/condition_evaluated
      -- 
    condition_evaluated_808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(19), ack => do_while_stmt_355_branch_req_0); -- 
    loadKernelChannel_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(86) & loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(23);
      gj_loadKernelChannel_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	24 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	23 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	43 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/aggregated_phi_sample_req
      -- CP-element group 20: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_sample_start__ps
      -- 
    loadKernelChannel_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(41) & loadKernelChannel_CP_671_elements(24) & loadKernelChannel_CP_671_elements(23);
      gj_loadKernelChannel_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	26 
    -- CP-element group 21: 	44 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	75 
    -- CP-element group 21: 	87 
    -- CP-element group 21: 	79 
    -- CP-element group 21: 	83 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	41 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/aggregated_phi_sample_ack
      -- CP-element group 21: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_sample_completed_
      -- 
    loadKernelChannel_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(26) & loadKernelChannel_CP_671_elements(44);
      gj_loadKernelChannel_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	42 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	45 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/aggregated_phi_update_req
      -- CP-element group 22: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_update_start__ps
      -- 
    loadKernelChannel_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(25) & loadKernelChannel_CP_671_elements(42);
      gj_loadKernelChannel_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	27 
    -- CP-element group 23: 	46 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/aggregated_phi_update_ack
      -- 
    loadKernelChannel_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(46);
      gj_loadKernelChannel_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	18 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	20 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_sample_start_
      -- 
    loadKernelChannel_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	18 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	72 
    -- CP-element group 25: 	27 
    -- CP-element group 25: 	61 
    -- CP-element group 25: 	66 
    -- CP-element group 25: 	80 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	22 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_update_start_
      -- 
    loadKernelChannel_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(72) & loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(66) & loadKernelChannel_CP_671_elements(80);
      gj_loadKernelChannel_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	70 
    -- CP-element group 27: 	78 
    -- CP-element group 27: 	60 
    -- CP-element group 27: 	66 
    -- CP-element group 27: 	19 
    -- CP-element group 27: 	23 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27:  members (15) 
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_resize_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_resize_1/index_resize_req
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_resized_1
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_resize_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_scale_1/$entry
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_resize_1/index_resize_ack
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_scale_1/$exit
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_scaled_1
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_computed_1
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_scale_1/scale_rename_req
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_index_scale_1/scale_rename_ack
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_update_completed__ps
      -- 
    req_960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(27), ack => array_obj_ref_402_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	16 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(28) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_loopback_sample_req
      -- CP-element group 29: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_loopback_sample_req_ps
      -- 
    phi_stmt_357_loopback_sample_req_823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_357_loopback_sample_req_823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(29), ack => phi_stmt_357_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(29) is bound as output of CP function.
    -- CP-element group 30:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(30) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 31:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_entry_sample_req
      -- CP-element group 31: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_entry_sample_req_ps
      -- 
    phi_stmt_357_entry_sample_req_826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_357_entry_sample_req_826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(31), ack => phi_stmt_357_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_phi_mux_ack
      -- CP-element group 32: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_357_phi_mux_ack_ps
      -- 
    phi_stmt_357_phi_mux_ack_829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_357_ack_0, ack => loadKernelChannel_CP_671_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_sample_start__ps
      -- CP-element group 33: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Sample/req
      -- 
    req_842_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_842_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(33), ack => nmycount_379_359_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_update_start__ps
      -- CP-element group 34: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_update_start_
      -- CP-element group 34: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Update/req
      -- 
    req_847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(34), ack => nmycount_379_359_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Sample/ack
      -- 
    ack_843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_379_359_buf_ack_0, ack => loadKernelChannel_CP_671_elements(35)); -- 
    -- CP-element group 36:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nmycount_359_Update/ack
      -- 
    ack_848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_379_359_buf_ack_1, ack => loadKernelChannel_CP_671_elements(36)); -- 
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_sample_start__ps
      -- CP-element group 37: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Sample/req
      -- 
    req_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(37), ack => start_add_360_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Update/req
      -- CP-element group 38: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_update_start__ps
      -- CP-element group 38: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_update_start_
      -- CP-element group 38: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Update/$entry
      -- 
    req_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(38), ack => start_add_360_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_sample_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Sample/ack
      -- 
    ack_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_360_buf_ack_0, ack => loadKernelChannel_CP_671_elements(39)); -- 
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_update_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_start_add_360_Update/$exit
      -- 
    ack_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_360_buf_ack_1, ack => loadKernelChannel_CP_671_elements(40)); -- 
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	18 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	77 
    -- CP-element group 41: 	85 
    -- CP-element group 41: 	81 
    -- CP-element group 41: 	21 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	20 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_sample_start_
      -- 
    loadKernelChannel_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(77) & loadKernelChannel_CP_671_elements(85) & loadKernelChannel_CP_671_elements(81) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	18 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	46 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	84 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	22 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_update_start_
      -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(61) & loadKernelChannel_CP_671_elements(84);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	20 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_sample_start__ps
      -- 
    loadKernelChannel_CP_671_elements(43) <= loadKernelChannel_CP_671_elements(20);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	21 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_sample_completed__ps
      -- 
    -- Element group loadKernelChannel_CP_671_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	22 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_update_start__ps
      -- 
    loadKernelChannel_CP_671_elements(45) <= loadKernelChannel_CP_671_elements(22);
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	60 
    -- CP-element group 46: 	82 
    -- CP-element group 46: 	23 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	42 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_update_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_update_completed_
      -- 
    -- Element group loadKernelChannel_CP_671_elements(46) is bound as output of CP function.
    -- CP-element group 47:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	16 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_loopback_trigger
      -- 
    loadKernelChannel_CP_671_elements(47) <= loadKernelChannel_CP_671_elements(16);
    -- CP-element group 48:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_loopback_sample_req
      -- CP-element group 48: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_loopback_sample_req_ps
      -- 
    phi_stmt_361_loopback_sample_req_877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_361_loopback_sample_req_877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(48), ack => phi_stmt_361_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(48) is bound as output of CP function.
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_entry_trigger
      -- 
    loadKernelChannel_CP_671_elements(49) <= loadKernelChannel_CP_671_elements(17);
    -- CP-element group 50:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_entry_sample_req
      -- CP-element group 50: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_entry_sample_req_ps
      -- 
    phi_stmt_361_entry_sample_req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_361_entry_sample_req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(50), ack => phi_stmt_361_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_phi_mux_ack
      -- CP-element group 51: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/phi_stmt_361_phi_mux_ack_ps
      -- 
    phi_stmt_361_phi_mux_ack_883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_361_ack_0, ack => loadKernelChannel_CP_671_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_sample_start__ps
      -- CP-element group 52: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Sample/req
      -- 
    req_896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(52), ack => nfetch_val_424_363_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_update_start__ps
      -- CP-element group 53: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_update_start_
      -- CP-element group 53: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Update/req
      -- 
    req_901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(53), ack => nfetch_val_424_363_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_sample_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Sample/$exit
      -- 
    ack_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_424_363_buf_ack_0, ack => loadKernelChannel_CP_671_elements(54)); -- 
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_update_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_nfetch_val_363_Update/ack
      -- 
    ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nfetch_val_424_363_buf_ack_1, ack => loadKernelChannel_CP_671_elements(55)); -- 
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_sample_start__ps
      -- CP-element group 56: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_sample_start_
      -- 
    req_914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(56), ack => my_fetch_344_364_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_671_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Update/req
      -- CP-element group 57: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_update_start__ps
      -- CP-element group 57: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_update_start_
      -- 
    req_919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(57), ack => my_fetch_344_364_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_671_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_sample_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_sample_completed_
      -- 
    ack_915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_344_364_buf_ack_0, ack => loadKernelChannel_CP_671_elements(58)); -- 
    -- CP-element group 59:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/R_my_fetch_364_update_completed__ps
      -- 
    ack_920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_fetch_344_364_buf_ack_1, ack => loadKernelChannel_CP_671_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	27 
    -- CP-element group 60: 	46 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Sample/req
      -- 
    req_929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(60), ack => WPIPE_kernel_pipe1_386_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	25 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_update_start_
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Update/req
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Sample/$exit
      -- 
    ack_930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_386_inst_ack_0, ack => loadKernelChannel_CP_671_elements(61)); -- 
    req_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(61), ack => WPIPE_kernel_pipe1_386_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	87 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Update/ack
      -- CP-element group 62: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/WPIPE_kernel_pipe1_386_Update/$exit
      -- 
    ack_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_386_inst_ack_1, ack => loadKernelChannel_CP_671_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	67 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	68 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_request/$entry
      -- CP-element group 63: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_request/req
      -- CP-element group 63: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_sample_start_
      -- 
    req_975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(63), ack => addr_of_403_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(67) & loadKernelChannel_CP_671_elements(68);
      gj_loadKernelChannel_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	18 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	76 
    -- CP-element group 64: 	69 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	69 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_complete/req
      -- CP-element group 64: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_update_start_
      -- 
    req_980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(64), ack => addr_of_403_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(76) & loadKernelChannel_CP_671_elements(69);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Update/req
      -- 
    req_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(65), ack => array_obj_ref_402_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(18) & loadKernelChannel_CP_671_elements(67) & loadKernelChannel_CP_671_elements(68);
      gj_loadKernelChannel_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	27 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	87 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	25 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_sample_complete
      -- CP-element group 66: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Sample/ack
      -- 
    ack_961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_index_offset_ack_0, ack => loadKernelChannel_CP_671_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	63 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (8) 
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_base_plus_offset/$entry
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_base_plus_offset/$exit
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_base_plus_offset/sum_rename_req
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_base_plus_offset/sum_rename_ack
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_root_address_calculated
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_offset_calculated
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/array_obj_ref_402_final_index_sum_regn_Update/ack
      -- 
    ack_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_index_offset_ack_1, ack => loadKernelChannel_CP_671_elements(67)); -- 
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	63 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: 	63 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_request/$exit
      -- CP-element group 68: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_request/ack
      -- CP-element group 68: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_sample_completed_
      -- 
    ack_976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_403_final_reg_ack_0, ack => loadKernelChannel_CP_671_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	64 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	64 
    -- CP-element group 69:  members (19) 
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_word_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_plus_offset/$exit
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_plus_offset/sum_rename_req
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_word_addrgen/$exit
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_word_addrgen/$entry
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_complete/$exit
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_plus_offset/sum_rename_ack
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_address_resized
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/addr_of_403_complete/ack
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_addr_resize/$exit
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_root_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_word_addrgen/root_register_req
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_addr_resize/base_resize_ack
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_plus_offset/$entry
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_addr_resize/$entry
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_address_calculated
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_base_addr_resize/base_resize_req
      -- CP-element group 69: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_word_addrgen/root_register_ack
      -- 
    ack_981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_403_final_reg_ack_1, ack => loadKernelChannel_CP_671_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	27 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Sample/req
      -- 
    req_989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(70), ack => W_fn_393_delayed_7_0_405_inst_req_0); -- 
    loadKernelChannel_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(72);
      gj_loadKernelChannel_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_update_start_
      -- CP-element group 71: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Update/req
      -- 
    req_994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(71), ack => W_fn_393_delayed_7_0_405_inst_req_1); -- 
    loadKernelChannel_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(73) & loadKernelChannel_CP_671_elements(76);
      gj_loadKernelChannel_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	25 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Sample/ack
      -- 
    ack_990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_393_delayed_7_0_405_inst_ack_0, ack => loadKernelChannel_CP_671_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_407_Update/ack
      -- 
    ack_995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_393_delayed_7_0_405_inst_ack_1, ack => loadKernelChannel_CP_671_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	69 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/word_0/rr
      -- CP-element group 74: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/word_0/$entry
      -- CP-element group 74: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/$entry
      -- CP-element group 74: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/$entry
      -- 
    rr_1028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(74), ack => ptr_deref_411_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(73) & loadKernelChannel_CP_671_elements(69) & loadKernelChannel_CP_671_elements(76);
      gj_loadKernelChannel_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	21 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/word_0/cr
      -- CP-element group 75: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/$entry
      -- CP-element group 75: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/word_0/$entry
      -- CP-element group 75: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_update_start_
      -- 
    cr_1039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(75), ack => ptr_deref_411_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(77);
      gj_loadKernelChannel_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	64 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/word_0/ra
      -- CP-element group 76: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/word_0/$exit
      -- CP-element group 76: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/word_access_start/$exit
      -- CP-element group 76: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_sample_completed_
      -- 
    ra_1029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_411_load_0_ack_0, ack => loadKernelChannel_CP_671_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	87 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	41 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/ptr_deref_411_Merge/$entry
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/ptr_deref_411_Merge/$exit
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/ptr_deref_411_Merge/merge_req
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/ptr_deref_411_Merge/merge_ack
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/word_0/ca
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/word_0/$exit
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_Update/word_access_complete/$exit
      -- CP-element group 77: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/ptr_deref_411_update_completed_
      -- 
    ca_1040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_411_load_0_ack_1, ack => loadKernelChannel_CP_671_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	27 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Sample/req
      -- 
    req_1053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(78), ack => W_fn_399_delayed_13_0_413_inst_req_0); -- 
    loadKernelChannel_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(27) & loadKernelChannel_CP_671_elements(80);
      gj_loadKernelChannel_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	21 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	81 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Update/req
      -- CP-element group 79: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_update_start_
      -- 
    req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1058_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(79), ack => W_fn_399_delayed_13_0_413_inst_req_1); -- 
    loadKernelChannel_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(81);
      gj_loadKernelChannel_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	25 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Sample/ack
      -- CP-element group 80: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_sample_completed_
      -- 
    ack_1054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_399_delayed_13_0_413_inst_ack_0, ack => loadKernelChannel_CP_671_elements(80)); -- 
    -- CP-element group 81:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	87 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	41 
    -- CP-element group 81: 	79 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_415_Update/ack
      -- 
    ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fn_399_delayed_13_0_413_inst_ack_1, ack => loadKernelChannel_CP_671_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	46 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Sample/req
      -- 
    req_1067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(82), ack => W_fetch_val_401_delayed_13_0_416_inst_req_0); -- 
    loadKernelChannel_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(46) & loadKernelChannel_CP_671_elements(84);
      gj_loadKernelChannel_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Update/req
      -- CP-element group 83: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_update_start_
      -- 
    req_1072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(83), ack => W_fetch_val_401_delayed_13_0_416_inst_req_1); -- 
    loadKernelChannel_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(21) & loadKernelChannel_CP_671_elements(85);
      gj_loadKernelChannel_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	42 
    -- CP-element group 84: 	82 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Sample/ack
      -- 
    ack_1068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_401_delayed_13_0_416_inst_ack_0, ack => loadKernelChannel_CP_671_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	41 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/assign_stmt_418_Update/ack
      -- 
    ack_1073_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_val_401_delayed_13_0_416_inst_ack_1, ack => loadKernelChannel_CP_671_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	18 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	19 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_671_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_671_elements(18), ack => loadKernelChannel_CP_671_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	77 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	62 
    -- CP-element group 87: 	66 
    -- CP-element group 87: 	81 
    -- CP-element group 87: 	21 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	15 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_354/do_while_stmt_355/do_while_stmt_355_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= loadKernelChannel_CP_671_elements(77) & loadKernelChannel_CP_671_elements(85) & loadKernelChannel_CP_671_elements(62) & loadKernelChannel_CP_671_elements(66) & loadKernelChannel_CP_671_elements(81) & loadKernelChannel_CP_671_elements(21);
      gj_loadKernelChannel_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_671_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	14 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_354/do_while_stmt_355/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_354/do_while_stmt_355/loop_exit/ack
      -- 
    ack_1078_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_355_branch_ack_0, ack => loadKernelChannel_CP_671_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	14 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_354/do_while_stmt_355/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_354/do_while_stmt_355/loop_taken/ack
      -- 
    ack_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_355_branch_ack_1, ack => loadKernelChannel_CP_671_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	12 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	10 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_354/do_while_stmt_355/$exit
      -- 
    loadKernelChannel_CP_671_elements(90) <= loadKernelChannel_CP_671_elements(12);
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	10 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 assign_stmt_438/type_cast_437_sample_completed_
      -- CP-element group 91: 	 assign_stmt_438/type_cast_437_Sample/$exit
      -- CP-element group 91: 	 assign_stmt_438/type_cast_437_Sample/ra
      -- 
    ra_1095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_437_inst_ack_0, ack => loadKernelChannel_CP_671_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	10 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 assign_stmt_438/type_cast_437_Update/ca
      -- CP-element group 92: 	 assign_stmt_438/WPIPE_size_pipe_433_Sample/$entry
      -- CP-element group 92: 	 assign_stmt_438/type_cast_437_Update/$exit
      -- CP-element group 92: 	 assign_stmt_438/WPIPE_size_pipe_433_Sample/req
      -- CP-element group 92: 	 assign_stmt_438/WPIPE_size_pipe_433_sample_start_
      -- CP-element group 92: 	 assign_stmt_438/type_cast_437_update_completed_
      -- 
    ca_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_437_inst_ack_1, ack => loadKernelChannel_CP_671_elements(92)); -- 
    req_1108_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1108_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(92), ack => WPIPE_size_pipe_433_inst_req_0); -- 
    -- CP-element group 93:  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (6) 
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_Update/$entry
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_Update/req
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_sample_completed_
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_Sample/ack
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_update_start_
      -- CP-element group 93: 	 assign_stmt_438/WPIPE_size_pipe_433_Sample/$exit
      -- 
    ack_1109_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_433_inst_ack_0, ack => loadKernelChannel_CP_671_elements(93)); -- 
    req_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_671_elements(93), ack => WPIPE_size_pipe_433_inst_req_1); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (5) 
      -- CP-element group 94: 	 assign_stmt_438/WPIPE_size_pipe_433_Update/ack
      -- CP-element group 94: 	 assign_stmt_438/$exit
      -- CP-element group 94: 	 assign_stmt_438/WPIPE_size_pipe_433_Update/$exit
      -- CP-element group 94: 	 $exit
      -- CP-element group 94: 	 assign_stmt_438/WPIPE_size_pipe_433_update_completed_
      -- 
    ack_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_433_inst_ack_1, ack => loadKernelChannel_CP_671_elements(94)); -- 
    loadKernelChannel_do_while_stmt_355_terminator_1083: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_355_terminator_1083", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_671_elements(15),loop_continue => loadKernelChannel_CP_671_elements(89),loop_terminate => loadKernelChannel_CP_671_elements(88),loop_back => loadKernelChannel_CP_671_elements(13),loop_exit => loadKernelChannel_CP_671_elements(12),clk => clk, reset => reset); -- 
    phi_stmt_357_phi_seq_867_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(28);
      loadKernelChannel_CP_671_elements(33)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(35);
      loadKernelChannel_CP_671_elements(34)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(36);
      loadKernelChannel_CP_671_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(30);
      loadKernelChannel_CP_671_elements(37)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(39);
      loadKernelChannel_CP_671_elements(38)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(40);
      loadKernelChannel_CP_671_elements(31) <= phi_mux_reqs(1);
      phi_stmt_357_phi_seq_867 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_357_phi_seq_867") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(20), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(26), 
          phi_update_req => loadKernelChannel_CP_671_elements(22), 
          phi_update_ack => loadKernelChannel_CP_671_elements(27), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(32), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_361_phi_seq_921_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_671_elements(47);
      loadKernelChannel_CP_671_elements(52)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_671_elements(54);
      loadKernelChannel_CP_671_elements(53)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_671_elements(55);
      loadKernelChannel_CP_671_elements(48) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_671_elements(49);
      loadKernelChannel_CP_671_elements(56)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_671_elements(58);
      loadKernelChannel_CP_671_elements(57)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_671_elements(59);
      loadKernelChannel_CP_671_elements(50) <= phi_mux_reqs(1);
      phi_stmt_361_phi_seq_921 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_361_phi_seq_921") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_671_elements(43), 
          phi_sample_ack => loadKernelChannel_CP_671_elements(44), 
          phi_update_req => loadKernelChannel_CP_671_elements(45), 
          phi_update_ack => loadKernelChannel_CP_671_elements(46), 
          phi_mux_ack => loadKernelChannel_CP_671_elements(51), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_809_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_671_elements(16);
        preds(1)  <= loadKernelChannel_CP_671_elements(17);
        entry_tmerge_809 : transition_merge -- 
          generic map(name => " entry_tmerge_809")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_671_elements(18));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u64_u64_370_wire : std_logic_vector(63 downto 0);
    signal AND_u64_u64_392_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_383_wire : std_logic_vector(63 downto 0);
    signal LSHR_u64_u64_401_resized : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_401_scaled : std_logic_vector(13 downto 0);
    signal LSHR_u64_u64_401_wire : std_logic_vector(63 downto 0);
    signal R_sh_start_337_resized : std_logic_vector(13 downto 0);
    signal R_sh_start_337_scaled : std_logic_vector(13 downto 0);
    signal SUB_u64_u64_371_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_429_wire : std_logic_vector(63 downto 0);
    signal SUB_u64_u64_436_wire : std_logic_vector(63 downto 0);
    signal ULT_u64_u1_430_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_338_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_338_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_338_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_338_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_338_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_338_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_402_root_address : std_logic_vector(13 downto 0);
    signal fetch_addr_340 : std_logic_vector(31 downto 0);
    signal fetch_addr_404 : std_logic_vector(31 downto 0);
    signal fetch_val_361 : std_logic_vector(63 downto 0);
    signal fetch_val_401_delayed_13_0_418 : std_logic_vector(63 downto 0);
    signal first_fill_349 : std_logic_vector(0 downto 0);
    signal fn_393_delayed_7_0_407 : std_logic_vector(0 downto 0);
    signal fn_395 : std_logic_vector(0 downto 0);
    signal fn_399_delayed_13_0_415 : std_logic_vector(0 downto 0);
    signal fv_412 : std_logic_vector(63 downto 0);
    signal konst_331_wire_constant : std_logic_vector(63 downto 0);
    signal konst_347_wire_constant : std_logic_vector(63 downto 0);
    signal konst_367_wire_constant : std_logic_vector(63 downto 0);
    signal konst_369_wire_constant : std_logic_vector(63 downto 0);
    signal konst_372_wire_constant : std_logic_vector(63 downto 0);
    signal konst_377_wire_constant : std_logic_vector(63 downto 0);
    signal konst_391_wire_constant : std_logic_vector(63 downto 0);
    signal konst_393_wire_constant : std_logic_vector(63 downto 0);
    signal konst_400_wire_constant : std_logic_vector(63 downto 0);
    signal konst_428_wire_constant : std_logic_vector(63 downto 0);
    signal my_fetch_344 : std_logic_vector(63 downto 0);
    signal my_fetch_344_364_buffered : std_logic_vector(63 downto 0);
    signal my_num1_374 : std_logic_vector(63 downto 0);
    signal mycount_357 : std_logic_vector(63 downto 0);
    signal nfetch_val_424 : std_logic_vector(63 downto 0);
    signal nfetch_val_424_363_buffered : std_logic_vector(63 downto 0);
    signal nmycount_379 : std_logic_vector(63 downto 0);
    signal nmycount_379_359_buffered : std_logic_vector(63 downto 0);
    signal ptr_deref_343_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_343_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_343_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_343_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_343_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_411_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_411_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_411_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_411_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_411_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_start_333 : std_logic_vector(63 downto 0);
    signal start_add_360_buffered : std_logic_vector(63 downto 0);
    signal start_next_353 : std_logic_vector(0 downto 0);
    signal type_cast_437_wire : std_logic_vector(31 downto 0);
    signal var_val_385 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_338_constant_part_of_offset <= "00000000000000";
    array_obj_ref_338_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_338_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_338_resized_base_address <= "00000000000000";
    array_obj_ref_402_constant_part_of_offset <= "00000000000000";
    array_obj_ref_402_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_402_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_402_resized_base_address <= "00000000000000";
    konst_331_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_347_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_367_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_369_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_372_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000100";
    konst_377_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_391_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    konst_393_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_400_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    konst_428_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    ptr_deref_343_word_offset_0 <= "00000000000000";
    ptr_deref_411_word_offset_0 <= "00000000000000";
    phi_stmt_357: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_379_359_buffered & start_add_360_buffered;
      req <= phi_stmt_357_req_0 & phi_stmt_357_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_357",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_357_ack_0,
          idata => idata,
          odata => mycount_357,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_357
    phi_stmt_361: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nfetch_val_424_363_buffered & my_fetch_344_364_buffered;
      req <= phi_stmt_361_req_0 & phi_stmt_361_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_361",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_361_ack_0,
          idata => idata,
          odata => fetch_val_361,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_361
    -- flow-through select operator MUX_423_inst
    nfetch_val_424 <= fv_412 when (fn_399_delayed_13_0_415(0) /=  '0') else fetch_val_401_delayed_13_0_418;
    W_fetch_val_401_delayed_13_0_416_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_val_401_delayed_13_0_416_inst_req_0;
      W_fetch_val_401_delayed_13_0_416_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_val_401_delayed_13_0_416_inst_req_1;
      W_fetch_val_401_delayed_13_0_416_inst_ack_1<= rack(0);
      W_fetch_val_401_delayed_13_0_416_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_val_401_delayed_13_0_416_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_val_361,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_val_401_delayed_13_0_418,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_393_delayed_7_0_405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_393_delayed_7_0_405_inst_req_0;
      W_fn_393_delayed_7_0_405_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_393_delayed_7_0_405_inst_req_1;
      W_fn_393_delayed_7_0_405_inst_ack_1<= rack(0);
      W_fn_393_delayed_7_0_405_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_393_delayed_7_0_405_inst",
        buffer_size => 7,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_393_delayed_7_0_407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fn_399_delayed_13_0_413_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fn_399_delayed_13_0_413_inst_req_0;
      W_fn_399_delayed_13_0_413_inst_ack_0<= wack(0);
      rreq(0) <= W_fn_399_delayed_13_0_413_inst_req_1;
      W_fn_399_delayed_13_0_413_inst_ack_1<= rack(0);
      W_fn_399_delayed_13_0_413_inst : InterlockBuffer generic map ( -- 
        name => "W_fn_399_delayed_13_0_413_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fn_395,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fn_399_delayed_13_0_415,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_339_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_339_final_reg_req_0;
      addr_of_339_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_339_final_reg_req_1;
      addr_of_339_final_reg_ack_1<= rack(0);
      addr_of_339_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_339_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_338_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_340,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_403_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_403_final_reg_req_0;
      addr_of_403_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_403_final_reg_req_1;
      addr_of_403_final_reg_ack_1<= rack(0);
      addr_of_403_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_403_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_402_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_404,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    my_fetch_344_364_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= my_fetch_344_364_buf_req_0;
      my_fetch_344_364_buf_ack_0<= wack(0);
      rreq(0) <= my_fetch_344_364_buf_req_1;
      my_fetch_344_364_buf_ack_1<= rack(0);
      my_fetch_344_364_buf : InterlockBuffer generic map ( -- 
        name => "my_fetch_344_364_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => my_fetch_344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => my_fetch_344_364_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nfetch_val_424_363_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nfetch_val_424_363_buf_req_0;
      nfetch_val_424_363_buf_ack_0<= wack(0);
      rreq(0) <= nfetch_val_424_363_buf_req_1;
      nfetch_val_424_363_buf_ack_1<= rack(0);
      nfetch_val_424_363_buf : InterlockBuffer generic map ( -- 
        name => "nfetch_val_424_363_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nfetch_val_424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nfetch_val_424_363_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_379_359_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_379_359_buf_req_0;
      nmycount_379_359_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_379_359_buf_req_1;
      nmycount_379_359_buf_ack_1<= rack(0);
      nmycount_379_359_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_379_359_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_379,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_379_359_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_360_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_360_buf_req_0;
      start_add_360_buf_ack_0<= wack(0);
      rreq(0) <= start_add_360_buf_req_1;
      start_add_360_buf_ack_1<= rack(0);
      start_add_360_buf : InterlockBuffer generic map ( -- 
        name => "start_add_360_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_360_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_384_inst
    process(LSHR_u64_u64_383_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := LSHR_u64_u64_383_wire(15 downto 0);
      var_val_385 <= tmp_var; -- 
    end process;
    type_cast_437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_437_inst_req_0;
      type_cast_437_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_437_inst_req_1;
      type_cast_437_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  first_fill_349(0);
      type_cast_437_inst_gI: SplitGuardInterface generic map(name => "type_cast_437_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => SUB_u64_u64_436_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_437_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_338_index_1_rename
    process(R_sh_start_337_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_sh_start_337_resized;
      ov(13 downto 0) := iv;
      R_sh_start_337_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_338_index_1_resize
    process(sh_start_333) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := sh_start_333;
      ov := iv(13 downto 0);
      R_sh_start_337_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_338_root_address_inst
    process(array_obj_ref_338_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_338_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_338_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_402_index_1_rename
    process(LSHR_u64_u64_401_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_401_resized;
      ov(13 downto 0) := iv;
      LSHR_u64_u64_401_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_402_index_1_resize
    process(LSHR_u64_u64_401_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LSHR_u64_u64_401_wire;
      ov := iv(13 downto 0);
      LSHR_u64_u64_401_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_402_root_address_inst
    process(array_obj_ref_402_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_402_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_402_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_addr_0
    process(ptr_deref_343_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_343_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_base_resize
    process(fetch_addr_340) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_340;
      ov := iv(13 downto 0);
      ptr_deref_343_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_gather_scatter
    process(ptr_deref_343_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_data_0;
      ov(63 downto 0) := iv;
      my_fetch_344 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_343_root_address_inst
    process(ptr_deref_343_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_343_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_343_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_411_addr_0
    process(ptr_deref_411_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_411_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_411_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_411_base_resize
    process(fetch_addr_404) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_404;
      ov := iv(13 downto 0);
      ptr_deref_411_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_411_gather_scatter
    process(ptr_deref_411_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_411_data_0;
      ov(63 downto 0) := iv;
      fv_412 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_411_root_address_inst
    process(ptr_deref_411_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_411_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_411_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_355_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u64_u1_430_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_355_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_355_branch_req_0,
          ack0 => do_while_stmt_355_branch_ack_0,
          ack1 => do_while_stmt_355_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_378_inst
    process(mycount_357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_357, konst_377_wire_constant, tmp_var);
      nmycount_379 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_370_inst
    process(mycount_357) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mycount_357, konst_369_wire_constant, tmp_var);
      AND_u64_u64_370_wire <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_392_inst
    process(nmycount_379) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(nmycount_379, konst_391_wire_constant, tmp_var);
      AND_u64_u64_392_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_348_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_347_wire_constant, tmp_var);
      first_fill_349 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_394_inst
    process(AND_u64_u64_392_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(AND_u64_u64_392_wire, konst_393_wire_constant, tmp_var);
      fn_395 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_332_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(start_add_buffer, konst_331_wire_constant, tmp_var);
      sh_start_333 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_383_inst
    process(fetch_val_361, my_num1_374) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(fetch_val_361, my_num1_374, tmp_var);
      LSHR_u64_u64_383_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_401_inst
    process(nmycount_379) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(nmycount_379, konst_400_wire_constant, tmp_var);
      LSHR_u64_u64_401_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_373_inst
    process(SUB_u64_u64_371_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(SUB_u64_u64_371_wire, konst_372_wire_constant, tmp_var);
      my_num1_374 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_371_inst
    process(konst_367_wire_constant, AND_u64_u64_370_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(konst_367_wire_constant, AND_u64_u64_370_wire, tmp_var);
      SUB_u64_u64_371_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_429_inst
    process(end_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, konst_428_wire_constant, tmp_var);
      SUB_u64_u64_429_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_436_inst
    process(end_add_buffer, start_add_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(end_add_buffer, start_add_buffer, tmp_var);
      SUB_u64_u64_436_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u64_u1_430_inst
    process(mycount_357, SUB_u64_u64_429_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_357, SUB_u64_u64_429_wire, tmp_var);
      ULT_u64_u1_430_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : array_obj_ref_338_index_offset 
    ApIntAdd_group_13: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_sh_start_337_scaled;
      array_obj_ref_338_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_338_index_offset_req_0;
      array_obj_ref_338_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_338_index_offset_req_1;
      array_obj_ref_338_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_13_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_402_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= LSHR_u64_u64_401_scaled;
      array_obj_ref_402_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_402_index_offset_req_0;
      array_obj_ref_402_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_402_index_offset_req_1;
      array_obj_ref_402_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_343_load_0 ptr_deref_411_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_343_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_411_load_0_req_0;
      ptr_deref_343_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_411_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_343_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_411_load_0_req_1;
      ptr_deref_343_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_411_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= fn_393_delayed_7_0_407(0);
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_343_word_address_0 & ptr_deref_411_word_address_0;
      ptr_deref_343_data_0 <= data_out(127 downto 64);
      ptr_deref_411_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_352_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_352_inst_req_0;
      RPIPE_input_done_pipe_352_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_352_inst_req_1;
      RPIPE_input_done_pipe_352_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_349(0);
      start_next_353 <= data_out(0 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_386_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_386_inst_req_0;
      WPIPE_kernel_pipe1_386_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_386_inst_req_1;
      WPIPE_kernel_pipe1_386_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= var_val_385;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_size_pipe_433_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_433_inst_req_0;
      WPIPE_size_pipe_433_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_433_inst_req_1;
      WPIPE_size_pipe_433_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= first_fill_349(0);
      data_in <= type_cast_437_wire;
      size_pipe_write_1_gI: SplitGuardInterface generic map(name => "size_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_637_start: Boolean;
  signal timer_CP_637_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_req_318_inst_req_0 : boolean;
  signal WPIPE_timer_req_318_inst_ack_0 : boolean;
  signal WPIPE_timer_req_318_inst_req_1 : boolean;
  signal WPIPE_timer_req_318_inst_ack_1 : boolean;
  signal RPIPE_timer_resp_323_inst_req_0 : boolean;
  signal RPIPE_timer_resp_323_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_323_inst_req_1 : boolean;
  signal RPIPE_timer_resp_323_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_637_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_637_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_637: Block -- control-path 
    signal timer_CP_637_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_637_elements(0) <= timer_CP_637_start;
    timer_CP_637_symbol <= timer_CP_637_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_sample_start_
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/req
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_sample_start_
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/rr
      -- 
    rr_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => RPIPE_timer_resp_323_inst_req_0); -- 
    req_650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(0), ack => WPIPE_timer_req_318_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_sample_completed_
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_update_start_
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Sample/ack
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/$entry
      -- CP-element group 1: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/req
      -- 
    ack_651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_318_inst_ack_0, ack => timer_CP_637_elements(1)); -- 
    req_655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(1), ack => WPIPE_timer_req_318_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_update_completed_
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/$exit
      -- CP-element group 2: 	 assign_stmt_321_to_assign_stmt_324/WPIPE_timer_req_318_Update/ack
      -- 
    ack_656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_318_inst_ack_1, ack => timer_CP_637_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_sample_completed_
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_update_start_
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Sample/ra
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/$entry
      -- CP-element group 3: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/cr
      -- 
    ra_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_323_inst_ack_0, ack => timer_CP_637_elements(3)); -- 
    cr_669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_637_elements(3), ack => RPIPE_timer_resp_323_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_update_completed_
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/$exit
      -- CP-element group 4: 	 assign_stmt_321_to_assign_stmt_324/RPIPE_timer_resp_323_Update/ca
      -- 
    ca_670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_323_inst_ack_1, ack => timer_CP_637_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_321_to_assign_stmt_324/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_637_elements(4) & timer_CP_637_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_637_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_320_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_320_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_323_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_323_inst_req_0;
      RPIPE_timer_resp_323_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_323_inst_req_1;
      RPIPE_timer_resp_323_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_318_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_318_inst_req_0;
      WPIPE_timer_req_318_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_318_inst_req_1;
      WPIPE_timer_req_318_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_320_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_4781_start: Boolean;
  signal timerDaemon_CP_4781_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_2104_req_1 : boolean;
  signal RPIPE_timer_req_2111_inst_ack_0 : boolean;
  signal RPIPE_timer_req_2111_inst_ack_1 : boolean;
  signal RPIPE_timer_req_2111_inst_req_0 : boolean;
  signal RPIPE_timer_req_2111_inst_req_1 : boolean;
  signal do_while_stmt_2102_branch_req_0 : boolean;
  signal phi_stmt_2104_req_0 : boolean;
  signal nCOUNTER_2117_2108_buf_ack_1 : boolean;
  signal nCOUNTER_2117_2108_buf_req_0 : boolean;
  signal nCOUNTER_2117_2108_buf_req_1 : boolean;
  signal nCOUNTER_2117_2108_buf_ack_0 : boolean;
  signal phi_stmt_2104_ack_0 : boolean;
  signal WPIPE_timer_resp_2119_inst_req_0 : boolean;
  signal WPIPE_timer_resp_2119_inst_ack_0 : boolean;
  signal WPIPE_timer_resp_2119_inst_req_1 : boolean;
  signal WPIPE_timer_resp_2119_inst_ack_1 : boolean;
  signal do_while_stmt_2102_branch_ack_0 : boolean;
  signal do_while_stmt_2102_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_4781_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4781_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_4781_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_4781_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_4781: Block -- control-path 
    signal timerDaemon_CP_4781_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_4781_elements(0) <= timerDaemon_CP_4781_start;
    timerDaemon_CP_4781_symbol <= timerDaemon_CP_4781_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_2101/do_while_stmt_2102__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2101/$entry
      -- CP-element group 0: 	 branch_block_stmt_2101/branch_block_stmt_2101__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_2101/do_while_stmt_2102__exit__
      -- CP-element group 1: 	 branch_block_stmt_2101/$exit
      -- CP-element group 1: 	 branch_block_stmt_2101/branch_block_stmt_2101__exit__
      -- CP-element group 1: 	 $exit
      -- 
    timerDaemon_CP_4781_elements(1) <= timerDaemon_CP_4781_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102__entry__
      -- CP-element group 2: 	 branch_block_stmt_2101/do_while_stmt_2102/$entry
      -- 
    timerDaemon_CP_4781_elements(2) <= timerDaemon_CP_4781_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102__exit__
      -- 
    -- Element group timerDaemon_CP_4781_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_back
      -- 
    -- Element group timerDaemon_CP_4781_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/$entry
      -- 
    timerDaemon_CP_4781_elements(5) <= timerDaemon_CP_4781_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_body_done
      -- 
    timerDaemon_CP_4781_elements(6) <= timerDaemon_CP_4781_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_4781_elements(7) <= timerDaemon_CP_4781_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_4781_elements(8) <= timerDaemon_CP_4781_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2109_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/loop_body_start
      -- 
    -- Element group timerDaemon_CP_4781_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/condition_evaluated
      -- 
    condition_evaluated_4805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(10), ack => do_while_stmt_2102_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(40) & timerDaemon_CP_4781_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: 	15 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(9) & timerDaemon_CP_4781_elements(15) & timerDaemon_CP_4781_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2109_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(35) & timerDaemon_CP_4781_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_update_req
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(32) & timerDaemon_CP_4781_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(36) & timerDaemon_CP_4781_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(9) & timerDaemon_CP_4781_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(9) & timerDaemon_CP_4781_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_4781_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_update_completed_
      -- 
    -- Element group timerDaemon_CP_4781_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_trigger
      -- 
    timerDaemon_CP_4781_elements(19) <= timerDaemon_CP_4781_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_loopback_sample_req_ps
      -- 
    phi_stmt_2104_loopback_sample_req_4820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2104_loopback_sample_req_4820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(20), ack => phi_stmt_2104_req_1); -- 
    -- Element group timerDaemon_CP_4781_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_trigger
      -- 
    timerDaemon_CP_4781_elements(21) <= timerDaemon_CP_4781_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_entry_sample_req
      -- 
    phi_stmt_2104_entry_sample_req_4823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2104_entry_sample_req_4823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(22), ack => phi_stmt_2104_req_0); -- 
    -- Element group timerDaemon_CP_4781_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2104_phi_mux_ack
      -- 
    phi_stmt_2104_phi_mux_ack_4826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2104_ack_0, ack => timerDaemon_CP_4781_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_sample_completed_
      -- 
    -- Element group timerDaemon_CP_4781_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_start_
      -- 
    -- Element group timerDaemon_CP_4781_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_completed__ps
      -- 
    timerDaemon_CP_4781_elements(26) <= timerDaemon_CP_4781_elements(27);
    -- CP-element group 27:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/type_cast_2107_update_completed_
      -- 
    -- Element group timerDaemon_CP_4781_elements(27) is a control-delay.
    cp_element_27_delay: control_delay_element  generic map(name => " 27_delay", delay_value => 1)  port map(req => timerDaemon_CP_4781_elements(25), ack => timerDaemon_CP_4781_elements(27), clk => clk, reset =>reset);
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Sample/req
      -- CP-element group 28: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Sample/$entry
      -- 
    req_4847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(28), ack => nCOUNTER_2117_2108_buf_req_0); -- 
    -- Element group timerDaemon_CP_4781_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_update_start_
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Update/req
      -- CP-element group 29: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_update_start__ps
      -- 
    req_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(29), ack => nCOUNTER_2117_2108_buf_req_1); -- 
    -- Element group timerDaemon_CP_4781_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Sample/ack
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_sample_completed_
      -- 
    ack_4848_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2117_2108_buf_ack_0, ack => timerDaemon_CP_4781_elements(30)); -- 
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/R_nCOUNTER_2108_update_completed__ps
      -- 
    ack_4853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_2117_2108_buf_ack_1, ack => timerDaemon_CP_4781_elements(31)); -- 
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2109_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(9) & timerDaemon_CP_4781_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Sample/$entry
      -- 
    rr_4866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(33), ack => RPIPE_timer_req_2111_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(11) & timerDaemon_CP_4781_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_update_start_
      -- CP-element group 34: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Update/cr
      -- 
    cr_4871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(34), ack => RPIPE_timer_req_2111_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(35) & timerDaemon_CP_4781_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_sample_completed_
      -- 
    ra_4867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2111_inst_ack_0, ack => timerDaemon_CP_4781_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/phi_stmt_2109_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/RPIPE_timer_req_2111_update_completed_
      -- 
    ca_4872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_2111_inst_ack_1, ack => timerDaemon_CP_4781_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Sample/req
      -- 
    req_4880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(37), ack => WPIPE_timer_resp_2119_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(36) & timerDaemon_CP_4781_elements(18) & timerDaemon_CP_4781_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_update_start_
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Update/req
      -- 
    ack_4881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2119_inst_ack_0, ack => timerDaemon_CP_4781_elements(38)); -- 
    req_4885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_4781_elements(38), ack => WPIPE_timer_resp_2119_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/WPIPE_timer_resp_2119_Update/ack
      -- 
    ack_4886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_2119_inst_ack_1, ack => timerDaemon_CP_4781_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_4781_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_4781_elements(9), ack => timerDaemon_CP_4781_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2101/do_while_stmt_2102/do_while_stmt_2102_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_4781_elements(39) & timerDaemon_CP_4781_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_4781_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_exit/ack
      -- 
    ack_4891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2102_branch_ack_0, ack => timerDaemon_CP_4781_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_2101/do_while_stmt_2102/loop_taken/ack
      -- 
    ack_4895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2102_branch_ack_1, ack => timerDaemon_CP_4781_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_2101/do_while_stmt_2102/$exit
      -- 
    timerDaemon_CP_4781_elements(44) <= timerDaemon_CP_4781_elements(3);
    timerDaemon_do_while_stmt_2102_terminator_4896: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_2102_terminator_4896", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_4781_elements(6),loop_continue => timerDaemon_CP_4781_elements(43),loop_terminate => timerDaemon_CP_4781_elements(42),loop_back => timerDaemon_CP_4781_elements(4),loop_exit => timerDaemon_CP_4781_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2104_phi_seq_4854_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_4781_elements(21);
      timerDaemon_CP_4781_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_4781_elements(24);
      timerDaemon_CP_4781_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_4781_elements(26);
      timerDaemon_CP_4781_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_4781_elements(19);
      timerDaemon_CP_4781_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_4781_elements(30);
      timerDaemon_CP_4781_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_4781_elements(31);
      timerDaemon_CP_4781_elements(20) <= phi_mux_reqs(1);
      phi_stmt_2104_phi_seq_4854 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_2104_phi_seq_4854") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_4781_elements(11), 
          phi_sample_ack => timerDaemon_CP_4781_elements(17), 
          phi_update_req => timerDaemon_CP_4781_elements(13), 
          phi_update_ack => timerDaemon_CP_4781_elements(18), 
          phi_mux_ack => timerDaemon_CP_4781_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4806_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_4781_elements(7);
        preds(1)  <= timerDaemon_CP_4781_elements(8);
        entry_tmerge_4806 : transition_merge -- 
          generic map(name => " entry_tmerge_4806")
          port map (preds => preds, symbol_out => timerDaemon_CP_4781_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_2104 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_2111_wire : std_logic_vector(0 downto 0);
    signal konst_2115_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2123_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_2117 : std_logic_vector(63 downto 0);
    signal nCOUNTER_2117_2108_buffered : std_logic_vector(63 downto 0);
    signal req_2109 : std_logic_vector(0 downto 0);
    signal type_cast_2107_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_2115_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_2123_wire_constant <= "1";
    type_cast_2107_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_2104: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2107_wire_constant & nCOUNTER_2117_2108_buffered;
      req <= phi_stmt_2104_req_0 & phi_stmt_2104_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2104",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2104_ack_0,
          idata => idata,
          odata => COUNTER_2104,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2104
    nCOUNTER_2117_2108_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_2117_2108_buf_req_0;
      nCOUNTER_2117_2108_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_2117_2108_buf_req_1;
      nCOUNTER_2117_2108_buf_ack_1<= rack(0);
      nCOUNTER_2117_2108_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_2117_2108_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_2117,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_2117_2108_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_2109
    process(RPIPE_timer_req_2111_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_2111_wire(0 downto 0);
      req_2109 <= tmp_var; -- 
    end process;
    do_while_stmt_2102_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2123_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2102_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2102_branch_req_0,
          ack0 => do_while_stmt_2102_branch_ack_0,
          ack1 => do_while_stmt_2102_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_2116_inst
    process(COUNTER_2104) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_2104, konst_2115_wire_constant, tmp_var);
      nCOUNTER_2117 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_2111_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_2111_inst_req_0;
      RPIPE_timer_req_2111_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_2111_inst_req_1;
      RPIPE_timer_req_2111_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_2111_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_2119_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_2119_inst_req_0;
      WPIPE_timer_resp_2119_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_2119_inst_req_1;
      WPIPE_timer_resp_2119_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_2109(0);
      data_in <= COUNTER_2104;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      num_cont : in  std_logic_vector(15 downto 0);
      row1 : in  std_logic_vector(15 downto 0);
      col1 : in  std_logic_vector(15 downto 0);
      rk1 : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_num_cont :  std_logic_vector(15 downto 0);
  signal access_T_row1 :  std_logic_vector(15 downto 0);
  signal access_T_col1 :  std_logic_vector(15 downto 0);
  signal access_T_rk1 :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(95 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(95 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(95 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(127 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(15 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(63 downto 0);
      end_add : in  std_logic_vector(63 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(15 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_end_add :  std_logic_vector(63 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(127 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(127 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(31 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(1 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(15 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_num_cont <= access_T_in_args(95 downto 80);
  access_T_row1 <= access_T_in_args(79 downto 64);
  access_T_col1 <= access_T_in_args(63 downto 48);
  access_T_rk1 <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 96,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      num_cont => access_T_num_cont,
      row1 => access_T_row1,
      col1 => access_T_col1,
      rk1 => access_T_rk1,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(15 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(95 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(127 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(15 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(15 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(0 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(15 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(127 downto 64);
  loadKernelChannel_end_add <= loadKernelChannel_in_args(63 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 128,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      end_add => loadKernelChannel_end_add,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(0 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(1 downto 1),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(1 downto 1),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(31 downto 16),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(31 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 100 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
