-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity access_T is -- 
  generic (tag_length : integer); 
  port ( -- 
    row_in : in  std_logic_vector(15 downto 0);
    chl_in : in  std_logic_vector(15 downto 0);
    ct : in  std_logic_vector(15 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
    input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
    input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
    input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity access_T;
architecture access_T_arch of access_T is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal row_in_buffer :  std_logic_vector(15 downto 0);
  signal row_in_update_enable: Boolean;
  signal chl_in_buffer :  std_logic_vector(15 downto 0);
  signal chl_in_update_enable: Boolean;
  signal ct_buffer :  std_logic_vector(15 downto 0);
  signal ct_update_enable: Boolean;
  -- output port buffer signals
  signal access_T_CP_0_start: Boolean;
  signal access_T_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_269_index_offset_req_0 : boolean;
  signal array_obj_ref_269_index_offset_ack_0 : boolean;
  signal WPIPE_input_pipe2_256_inst_ack_1 : boolean;
  signal n_start4_344_123_buf_req_1 : boolean;
  signal n_row4_363_120_buf_req_1 : boolean;
  signal array_obj_ref_269_index_offset_req_1 : boolean;
  signal array_obj_ref_269_index_offset_ack_1 : boolean;
  signal n_row4_363_120_buf_ack_1 : boolean;
  signal phi_stmt_44_req_0 : boolean;
  signal addr_of_204_final_reg_ack_1 : boolean;
  signal addr_of_138_final_reg_req_1 : boolean;
  signal do_while_stmt_42_branch_req_0 : boolean;
  signal W_send_flag2_249_delayed_13_0_252_inst_ack_0 : boolean;
  signal addr_of_204_final_reg_req_1 : boolean;
  signal phi_stmt_44_req_1 : boolean;
  signal WPIPE_input_pipe2_256_inst_req_1 : boolean;
  signal n_row4_363_120_buf_ack_0 : boolean;
  signal phi_stmt_44_ack_0 : boolean;
  signal addr_of_138_final_reg_ack_0 : boolean;
  signal addr_of_138_final_reg_req_0 : boolean;
  signal ptr_deref_208_load_0_ack_0 : boolean;
  signal ptr_deref_208_load_0_req_0 : boolean;
  signal n_address1_175_48_buf_req_0 : boolean;
  signal n_address1_175_48_buf_ack_0 : boolean;
  signal n_row4_363_120_buf_req_0 : boolean;
  signal n_address1_175_48_buf_req_1 : boolean;
  signal n_address1_175_48_buf_ack_1 : boolean;
  signal array_obj_ref_203_index_offset_ack_1 : boolean;
  signal phi_stmt_49_req_1 : boolean;
  signal W_send_flag1_186_delayed_13_0_186_inst_ack_1 : boolean;
  signal phi_stmt_49_req_0 : boolean;
  signal W_send_flag1_186_delayed_13_0_186_inst_req_1 : boolean;
  signal phi_stmt_49_ack_0 : boolean;
  signal type_cast_52_inst_req_0 : boolean;
  signal type_cast_52_inst_ack_0 : boolean;
  signal type_cast_52_inst_req_1 : boolean;
  signal type_cast_52_inst_ack_1 : boolean;
  signal n_address2_241_66_buf_req_1 : boolean;
  signal n_address2_241_66_buf_ack_1 : boolean;
  signal n_mycounter1_157_53_buf_req_0 : boolean;
  signal n_mycounter1_157_53_buf_ack_0 : boolean;
  signal array_obj_ref_203_index_offset_req_1 : boolean;
  signal n_mycounter1_157_53_buf_req_1 : boolean;
  signal n_mycounter1_157_53_buf_ack_1 : boolean;
  signal n_start4_344_123_buf_ack_0 : boolean;
  signal n_start4_344_123_buf_req_0 : boolean;
  signal W_send_flag1_186_delayed_13_0_186_inst_ack_0 : boolean;
  signal W_send_flag1_186_delayed_13_0_186_inst_req_0 : boolean;
  signal phi_stmt_54_req_1 : boolean;
  signal phi_stmt_54_req_0 : boolean;
  signal phi_stmt_54_ack_0 : boolean;
  signal addr_of_204_final_reg_ack_0 : boolean;
  signal array_obj_ref_137_index_offset_ack_1 : boolean;
  signal W_send_flag2_249_delayed_13_0_252_inst_req_0 : boolean;
  signal array_obj_ref_137_index_offset_req_1 : boolean;
  signal n_row1_165_58_buf_req_0 : boolean;
  signal n_row1_165_58_buf_ack_0 : boolean;
  signal n_row1_165_58_buf_req_1 : boolean;
  signal n_row1_165_58_buf_ack_1 : boolean;
  signal array_obj_ref_137_index_offset_ack_0 : boolean;
  signal array_obj_ref_203_index_offset_ack_0 : boolean;
  signal array_obj_ref_203_index_offset_req_0 : boolean;
  signal phi_stmt_59_req_0 : boolean;
  signal phi_stmt_59_req_1 : boolean;
  signal phi_stmt_59_ack_0 : boolean;
  signal array_obj_ref_137_index_offset_req_0 : boolean;
  signal n_start1_146_61_buf_req_0 : boolean;
  signal n_start1_146_61_buf_ack_0 : boolean;
  signal W_send_flag2_249_delayed_13_0_252_inst_ack_1 : boolean;
  signal n_start1_146_61_buf_req_1 : boolean;
  signal n_start1_146_61_buf_ack_1 : boolean;
  signal addr_of_204_final_reg_req_0 : boolean;
  signal phi_stmt_64_req_0 : boolean;
  signal phi_stmt_64_req_1 : boolean;
  signal WPIPE_input_pipe2_256_inst_ack_0 : boolean;
  signal phi_stmt_64_ack_0 : boolean;
  signal n_address2_241_66_buf_req_0 : boolean;
  signal n_address2_241_66_buf_ack_0 : boolean;
  signal phi_stmt_94_req_1 : boolean;
  signal phi_stmt_94_req_0 : boolean;
  signal type_cast_68_inst_req_0 : boolean;
  signal type_cast_68_inst_ack_0 : boolean;
  signal type_cast_68_inst_req_1 : boolean;
  signal type_cast_68_inst_ack_1 : boolean;
  signal W_send_flag2_249_delayed_13_0_252_inst_req_1 : boolean;
  signal phi_stmt_69_req_0 : boolean;
  signal ptr_deref_142_load_0_ack_1 : boolean;
  signal phi_stmt_69_req_1 : boolean;
  signal ptr_deref_142_load_0_req_1 : boolean;
  signal WPIPE_input_pipe2_256_inst_req_0 : boolean;
  signal phi_stmt_69_ack_0 : boolean;
  signal n_mycounter2_223_71_buf_req_0 : boolean;
  signal n_mycounter2_223_71_buf_ack_0 : boolean;
  signal n_mycounter2_223_71_buf_req_1 : boolean;
  signal n_mycounter2_223_71_buf_ack_1 : boolean;
  signal type_cast_73_inst_req_0 : boolean;
  signal type_cast_73_inst_ack_0 : boolean;
  signal type_cast_73_inst_req_1 : boolean;
  signal type_cast_73_inst_ack_1 : boolean;
  signal n_start4_344_123_buf_ack_1 : boolean;
  signal phi_stmt_74_req_1 : boolean;
  signal phi_stmt_74_req_0 : boolean;
  signal ptr_deref_142_load_0_ack_0 : boolean;
  signal phi_stmt_74_ack_0 : boolean;
  signal ptr_deref_142_load_0_req_0 : boolean;
  signal n_row2_231_78_buf_req_0 : boolean;
  signal n_row2_231_78_buf_ack_0 : boolean;
  signal n_row2_231_78_buf_req_1 : boolean;
  signal n_row2_231_78_buf_ack_1 : boolean;
  signal addr_of_138_final_reg_ack_1 : boolean;
  signal phi_stmt_79_req_1 : boolean;
  signal phi_stmt_79_req_0 : boolean;
  signal ptr_deref_208_load_0_ack_1 : boolean;
  signal phi_stmt_79_ack_0 : boolean;
  signal WPIPE_input_pipe1_190_inst_ack_1 : boolean;
  signal WPIPE_input_pipe1_190_inst_req_1 : boolean;
  signal n_start2_212_83_buf_req_0 : boolean;
  signal n_start2_212_83_buf_ack_0 : boolean;
  signal n_start2_212_83_buf_req_1 : boolean;
  signal n_start2_212_83_buf_ack_1 : boolean;
  signal phi_stmt_121_ack_0 : boolean;
  signal phi_stmt_84_req_0 : boolean;
  signal phi_stmt_84_req_1 : boolean;
  signal ptr_deref_208_load_0_req_1 : boolean;
  signal phi_stmt_116_ack_0 : boolean;
  signal phi_stmt_84_ack_0 : boolean;
  signal n_address3_307_86_buf_req_0 : boolean;
  signal n_address3_307_86_buf_ack_0 : boolean;
  signal n_address3_307_86_buf_req_1 : boolean;
  signal n_address3_307_86_buf_ack_1 : boolean;
  signal type_cast_88_inst_req_0 : boolean;
  signal type_cast_88_inst_ack_0 : boolean;
  signal type_cast_88_inst_req_1 : boolean;
  signal type_cast_88_inst_ack_1 : boolean;
  signal phi_stmt_116_req_0 : boolean;
  signal phi_stmt_121_req_1 : boolean;
  signal WPIPE_input_pipe1_190_inst_ack_0 : boolean;
  signal WPIPE_input_pipe1_190_inst_req_0 : boolean;
  signal phi_stmt_89_req_0 : boolean;
  signal phi_stmt_89_req_1 : boolean;
  signal phi_stmt_89_ack_0 : boolean;
  signal phi_stmt_121_req_0 : boolean;
  signal n_mycounter3_289_91_buf_req_0 : boolean;
  signal n_mycounter3_289_91_buf_ack_0 : boolean;
  signal n_mycounter3_289_91_buf_req_1 : boolean;
  signal n_mycounter3_289_91_buf_ack_1 : boolean;
  signal phi_stmt_116_req_1 : boolean;
  signal type_cast_93_inst_req_0 : boolean;
  signal type_cast_93_inst_ack_0 : boolean;
  signal type_cast_93_inst_req_1 : boolean;
  signal type_cast_93_inst_ack_1 : boolean;
  signal phi_stmt_94_ack_0 : boolean;
  signal n_row3_297_98_buf_req_0 : boolean;
  signal n_row3_297_98_buf_ack_0 : boolean;
  signal n_row3_297_98_buf_req_1 : boolean;
  signal n_row3_297_98_buf_ack_1 : boolean;
  signal phi_stmt_99_req_0 : boolean;
  signal phi_stmt_99_req_1 : boolean;
  signal phi_stmt_99_ack_0 : boolean;
  signal n_start3_278_101_buf_req_0 : boolean;
  signal n_start3_278_101_buf_ack_0 : boolean;
  signal n_start3_278_101_buf_req_1 : boolean;
  signal n_start3_278_101_buf_ack_1 : boolean;
  signal phi_stmt_104_req_1 : boolean;
  signal phi_stmt_104_req_0 : boolean;
  signal phi_stmt_104_ack_0 : boolean;
  signal type_cast_109_inst_req_0 : boolean;
  signal type_cast_109_inst_ack_0 : boolean;
  signal type_cast_109_inst_req_1 : boolean;
  signal type_cast_109_inst_ack_1 : boolean;
  signal n_address4_373_110_buf_req_0 : boolean;
  signal n_address4_373_110_buf_ack_0 : boolean;
  signal n_address4_373_110_buf_req_1 : boolean;
  signal n_address4_373_110_buf_ack_1 : boolean;
  signal phi_stmt_111_req_0 : boolean;
  signal phi_stmt_111_req_1 : boolean;
  signal phi_stmt_111_ack_0 : boolean;
  signal n_mycounter4_355_113_buf_req_0 : boolean;
  signal n_mycounter4_355_113_buf_ack_0 : boolean;
  signal n_mycounter4_355_113_buf_req_1 : boolean;
  signal n_mycounter4_355_113_buf_ack_1 : boolean;
  signal type_cast_115_inst_req_0 : boolean;
  signal type_cast_115_inst_ack_0 : boolean;
  signal type_cast_115_inst_req_1 : boolean;
  signal type_cast_115_inst_ack_1 : boolean;
  signal addr_of_270_final_reg_req_0 : boolean;
  signal addr_of_270_final_reg_ack_0 : boolean;
  signal addr_of_270_final_reg_req_1 : boolean;
  signal addr_of_270_final_reg_ack_1 : boolean;
  signal ptr_deref_274_load_0_req_0 : boolean;
  signal ptr_deref_274_load_0_ack_0 : boolean;
  signal ptr_deref_274_load_0_req_1 : boolean;
  signal ptr_deref_274_load_0_ack_1 : boolean;
  signal W_send_flag3_312_delayed_13_0_318_inst_req_0 : boolean;
  signal W_send_flag3_312_delayed_13_0_318_inst_ack_0 : boolean;
  signal W_send_flag3_312_delayed_13_0_318_inst_req_1 : boolean;
  signal W_send_flag3_312_delayed_13_0_318_inst_ack_1 : boolean;
  signal WPIPE_input_pipe3_322_inst_req_0 : boolean;
  signal WPIPE_input_pipe3_322_inst_ack_0 : boolean;
  signal WPIPE_input_pipe3_322_inst_req_1 : boolean;
  signal WPIPE_input_pipe3_322_inst_ack_1 : boolean;
  signal array_obj_ref_335_index_offset_req_0 : boolean;
  signal array_obj_ref_335_index_offset_ack_0 : boolean;
  signal array_obj_ref_335_index_offset_req_1 : boolean;
  signal array_obj_ref_335_index_offset_ack_1 : boolean;
  signal addr_of_336_final_reg_req_0 : boolean;
  signal addr_of_336_final_reg_ack_0 : boolean;
  signal addr_of_336_final_reg_req_1 : boolean;
  signal addr_of_336_final_reg_ack_1 : boolean;
  signal ptr_deref_340_load_0_req_0 : boolean;
  signal ptr_deref_340_load_0_ack_0 : boolean;
  signal ptr_deref_340_load_0_req_1 : boolean;
  signal ptr_deref_340_load_0_ack_1 : boolean;
  signal W_send_flag4_375_delayed_13_0_384_inst_req_0 : boolean;
  signal W_send_flag4_375_delayed_13_0_384_inst_ack_0 : boolean;
  signal W_send_flag4_375_delayed_13_0_384_inst_req_1 : boolean;
  signal W_send_flag4_375_delayed_13_0_384_inst_ack_1 : boolean;
  signal WPIPE_input_pipe4_388_inst_req_0 : boolean;
  signal WPIPE_input_pipe4_388_inst_ack_0 : boolean;
  signal WPIPE_input_pipe4_388_inst_req_1 : boolean;
  signal WPIPE_input_pipe4_388_inst_ack_1 : boolean;
  signal do_while_stmt_42_branch_ack_0 : boolean;
  signal do_while_stmt_42_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "access_T_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(15 downto 0) <= row_in;
  row_in_buffer <= in_buffer_data_out(15 downto 0);
  in_buffer_data_in(31 downto 16) <= chl_in;
  chl_in_buffer <= in_buffer_data_out(31 downto 16);
  in_buffer_data_in(47 downto 32) <= ct;
  ct_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  access_T_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "access_T_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= access_T_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  access_T_CP_0: Block -- control-path 
    signal access_T_CP_0_elements: BooleanArray(407 downto 0);
    -- 
  begin -- 
    access_T_CP_0_elements(0) <= access_T_CP_0_start;
    access_T_CP_0_symbol <= access_T_CP_0_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41__exit__
      -- CP-element group 0: 	 branch_block_stmt_29/do_while_stmt_42__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_29/$entry
      -- CP-element group 0: 	 branch_block_stmt_29/branch_block_stmt_29__entry__
      -- CP-element group 0: 	 branch_block_stmt_29/assign_stmt_36_to_assign_stmt_41__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	407 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_29/do_while_stmt_42__exit__
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_29/$exit
      -- CP-element group 1: 	 branch_block_stmt_29/branch_block_stmt_29__exit__
      -- 
    access_T_CP_0_elements(1) <= access_T_CP_0_elements(407);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_29/do_while_stmt_42/$entry
      -- CP-element group 2: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42__entry__
      -- 
    access_T_CP_0_elements(2) <= access_T_CP_0_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	407 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42__exit__
      -- 
    -- Element group access_T_CP_0_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_29/do_while_stmt_42/loop_back
      -- 
    -- Element group access_T_CP_0_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	405 
    -- CP-element group 5: 	406 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/condition_done
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/$entry
      -- 
    access_T_CP_0_elements(5) <= access_T_CP_0_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	404 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_29/do_while_stmt_42/loop_body_done
      -- 
    access_T_CP_0_elements(6) <= access_T_CP_0_elements(404);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	318 
    -- CP-element group 7: 	200 
    -- CP-element group 7: 	240 
    -- CP-element group 7: 	221 
    -- CP-element group 7: 	259 
    -- CP-element group 7: 	21 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	61 
    -- CP-element group 7: 	80 
    -- CP-element group 7: 	280 
    -- CP-element group 7: 	301 
    -- CP-element group 7: 	99 
    -- CP-element group 7: 	120 
    -- CP-element group 7: 	141 
    -- CP-element group 7: 	160 
    -- CP-element group 7: 	179 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/back_edge_to_loop_body
      -- 
    access_T_CP_0_elements(7) <= access_T_CP_0_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	242 
    -- CP-element group 8: 	202 
    -- CP-element group 8: 	223 
    -- CP-element group 8: 	261 
    -- CP-element group 8: 	23 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	63 
    -- CP-element group 8: 	82 
    -- CP-element group 8: 	282 
    -- CP-element group 8: 	303 
    -- CP-element group 8: 	320 
    -- CP-element group 8: 	101 
    -- CP-element group 8: 	122 
    -- CP-element group 8: 	143 
    -- CP-element group 8: 	162 
    -- CP-element group 8: 	181 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/first_time_through_loop_body
      -- 
    access_T_CP_0_elements(8) <= access_T_CP_0_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	314 
    -- CP-element group 9: 	315 
    -- CP-element group 9: 	195 
    -- CP-element group 9: 	234 
    -- CP-element group 9: 	194 
    -- CP-element group 9: 	216 
    -- CP-element group 9: 	235 
    -- CP-element group 9: 	215 
    -- CP-element group 9: 	254 
    -- CP-element group 9: 	253 
    -- CP-element group 9: 	333 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	56 
    -- CP-element group 9: 	74 
    -- CP-element group 9: 	75 
    -- CP-element group 9: 	368 
    -- CP-element group 9: 	369 
    -- CP-element group 9: 	386 
    -- CP-element group 9: 	387 
    -- CP-element group 9: 	403 
    -- CP-element group 9: 	274 
    -- CP-element group 9: 	275 
    -- CP-element group 9: 	295 
    -- CP-element group 9: 	296 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	332 
    -- CP-element group 9: 	350 
    -- CP-element group 9: 	351 
    -- CP-element group 9: 	93 
    -- CP-element group 9: 	94 
    -- CP-element group 9: 	114 
    -- CP-element group 9: 	115 
    -- CP-element group 9: 	135 
    -- CP-element group 9: 	136 
    -- CP-element group 9: 	154 
    -- CP-element group 9: 	155 
    -- CP-element group 9: 	173 
    -- CP-element group 9: 	174 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/loop_body_start
      -- 
    -- Element group access_T_CP_0_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	403 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/condition_evaluated
      -- 
    condition_evaluated_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(10), ack => do_while_stmt_42_branch_req_0); -- 
    access_T_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(403) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	314 
    -- CP-element group 11: 	234 
    -- CP-element group 11: 	194 
    -- CP-element group 11: 	215 
    -- CP-element group 11: 	253 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	55 
    -- CP-element group 11: 	74 
    -- CP-element group 11: 	274 
    -- CP-element group 11: 	295 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	93 
    -- CP-element group 11: 	114 
    -- CP-element group 11: 	135 
    -- CP-element group 11: 	154 
    -- CP-element group 11: 	173 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	255 
    -- CP-element group 11: 	217 
    -- CP-element group 11: 	236 
    -- CP-element group 11: 	196 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	57 
    -- CP-element group 11: 	76 
    -- CP-element group 11: 	276 
    -- CP-element group 11: 	297 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	116 
    -- CP-element group 11: 	137 
    -- CP-element group 11: 	156 
    -- CP-element group 11: 	175 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_start__ps
      -- 
    access_T_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= access_T_CP_0_elements(314) & access_T_CP_0_elements(234) & access_T_CP_0_elements(194) & access_T_CP_0_elements(215) & access_T_CP_0_elements(253) & access_T_CP_0_elements(34) & access_T_CP_0_elements(55) & access_T_CP_0_elements(74) & access_T_CP_0_elements(274) & access_T_CP_0_elements(295) & access_T_CP_0_elements(15) & access_T_CP_0_elements(93) & access_T_CP_0_elements(114) & access_T_CP_0_elements(135) & access_T_CP_0_elements(154) & access_T_CP_0_elements(173) & access_T_CP_0_elements(14);
      gj_access_T_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	316 
    -- CP-element group 12: 	197 
    -- CP-element group 12: 	237 
    -- CP-element group 12: 	218 
    -- CP-element group 12: 	256 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	58 
    -- CP-element group 12: 	77 
    -- CP-element group 12: 	277 
    -- CP-element group 12: 	298 
    -- CP-element group 12: 	96 
    -- CP-element group 12: 	117 
    -- CP-element group 12: 	138 
    -- CP-element group 12: 	157 
    -- CP-element group 12: 	176 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	404 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	314 
    -- CP-element group 12: 	234 
    -- CP-element group 12: 	194 
    -- CP-element group 12: 	215 
    -- CP-element group 12: 	253 
    -- CP-element group 12: 	34 
    -- CP-element group 12: 	55 
    -- CP-element group 12: 	74 
    -- CP-element group 12: 	274 
    -- CP-element group 12: 	295 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	93 
    -- CP-element group 12: 	114 
    -- CP-element group 12: 	135 
    -- CP-element group 12: 	154 
    -- CP-element group 12: 	173 
    -- CP-element group 12:  members (17) 
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_completed_
      -- 
    access_T_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(316) & access_T_CP_0_elements(197) & access_T_CP_0_elements(237) & access_T_CP_0_elements(218) & access_T_CP_0_elements(256) & access_T_CP_0_elements(18) & access_T_CP_0_elements(37) & access_T_CP_0_elements(58) & access_T_CP_0_elements(77) & access_T_CP_0_elements(277) & access_T_CP_0_elements(298) & access_T_CP_0_elements(96) & access_T_CP_0_elements(117) & access_T_CP_0_elements(138) & access_T_CP_0_elements(157) & access_T_CP_0_elements(176);
      gj_access_T_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	315 
    -- CP-element group 13: 	195 
    -- CP-element group 13: 	216 
    -- CP-element group 13: 	235 
    -- CP-element group 13: 	254 
    -- CP-element group 13: 	35 
    -- CP-element group 13: 	56 
    -- CP-element group 13: 	75 
    -- CP-element group 13: 	275 
    -- CP-element group 13: 	296 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	94 
    -- CP-element group 13: 	115 
    -- CP-element group 13: 	136 
    -- CP-element group 13: 	155 
    -- CP-element group 13: 	174 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	198 
    -- CP-element group 13: 	238 
    -- CP-element group 13: 	219 
    -- CP-element group 13: 	257 
    -- CP-element group 13: 	19 
    -- CP-element group 13: 	38 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	78 
    -- CP-element group 13: 	278 
    -- CP-element group 13: 	299 
    -- CP-element group 13: 	97 
    -- CP-element group 13: 	118 
    -- CP-element group 13: 	139 
    -- CP-element group 13: 	158 
    -- CP-element group 13: 	177 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_start__ps
      -- 
    access_T_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(315) & access_T_CP_0_elements(195) & access_T_CP_0_elements(216) & access_T_CP_0_elements(235) & access_T_CP_0_elements(254) & access_T_CP_0_elements(35) & access_T_CP_0_elements(56) & access_T_CP_0_elements(75) & access_T_CP_0_elements(275) & access_T_CP_0_elements(296) & access_T_CP_0_elements(16) & access_T_CP_0_elements(94) & access_T_CP_0_elements(115) & access_T_CP_0_elements(136) & access_T_CP_0_elements(155) & access_T_CP_0_elements(174);
      gj_access_T_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	317 
    -- CP-element group 14: 	199 
    -- CP-element group 14: 	220 
    -- CP-element group 14: 	239 
    -- CP-element group 14: 	258 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	60 
    -- CP-element group 14: 	79 
    -- CP-element group 14: 	279 
    -- CP-element group 14: 	300 
    -- CP-element group 14: 	98 
    -- CP-element group 14: 	119 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	159 
    -- CP-element group 14: 	178 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/aggregated_phi_update_ack
      -- 
    access_T_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 15) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15,11 => 15,12 => 15,13 => 15,14 => 15,15 => 15);
      constant place_markings: IntegerArray(0 to 15)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant place_delays: IntegerArray(0 to 15) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 16); -- 
    begin -- 
      preds <= access_T_CP_0_elements(317) & access_T_CP_0_elements(199) & access_T_CP_0_elements(220) & access_T_CP_0_elements(239) & access_T_CP_0_elements(258) & access_T_CP_0_elements(20) & access_T_CP_0_elements(39) & access_T_CP_0_elements(60) & access_T_CP_0_elements(79) & access_T_CP_0_elements(279) & access_T_CP_0_elements(300) & access_T_CP_0_elements(98) & access_T_CP_0_elements(119) & access_T_CP_0_elements(140) & access_T_CP_0_elements(159) & access_T_CP_0_elements(178);
      gj_access_T_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 16, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_start_
      -- 
    access_T_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	334 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_start_
      -- 
    access_T_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(334);
      gj_access_T_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_start__ps
      -- 
    access_T_CP_0_elements(17) <= access_T_CP_0_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_start__ps
      -- 
    access_T_CP_0_elements(19) <= access_T_CP_0_elements(13);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	334 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (15) 
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_scale_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_scale_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Sample/req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_scale_1/scale_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_scale_1/scale_rename_req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_resize_1/index_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_resize_1/index_resize_req
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_resize_1/$exit
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_resize_1/$entry
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_computed_1
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_scaled_1
      -- CP-element group 20: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_index_resized_1
      -- 
    req_833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(20), ack => array_obj_ref_137_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_trigger
      -- 
    access_T_CP_0_elements(21) <= access_T_CP_0_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_loopback_sample_req_ps
      -- 
    phi_stmt_44_loopback_sample_req_44_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_44_loopback_sample_req_44_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(22), ack => phi_stmt_44_req_1); -- 
    -- Element group access_T_CP_0_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_trigger
      -- 
    access_T_CP_0_elements(23) <= access_T_CP_0_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_sample_req
      -- CP-element group 24: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_entry_sample_req_ps
      -- 
    phi_stmt_44_entry_sample_req_47_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_44_entry_sample_req_47_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(24), ack => phi_stmt_44_req_0); -- 
    -- Element group access_T_CP_0_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_44_phi_mux_ack_ps
      -- 
    phi_stmt_44_phi_mux_ack_50_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_44_ack_0, ack => access_T_CP_0_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_start_
      -- 
    -- Element group access_T_CP_0_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_completed__ps
      -- 
    access_T_CP_0_elements(28) <= access_T_CP_0_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_47_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(27), ack => access_T_CP_0_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_start__ps
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/req
      -- 
    req_71_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_71_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(30), ack => n_address1_175_48_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_start__ps
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_start_
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/req
      -- 
    req_76_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_76_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(31), ack => n_address1_175_48_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Sample/ack
      -- 
    ack_72_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_175_48_buf_ack_0, ack => access_T_CP_0_elements(32)); -- 
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address1_48_Update/ack
      -- 
    ack_77_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_175_48_buf_ack_1, ack => access_T_CP_0_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	12 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	11 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_start_
      -- 
    access_T_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	39 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	13 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_start_
      -- 
    access_T_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(39);
      gj_access_T_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_start__ps
      -- 
    access_T_CP_0_elements(36) <= access_T_CP_0_elements(11);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_start__ps
      -- 
    access_T_CP_0_elements(38) <= access_T_CP_0_elements(13);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	35 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_trigger
      -- 
    access_T_CP_0_elements(40) <= access_T_CP_0_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_loopback_sample_req_ps
      -- 
    phi_stmt_49_loopback_sample_req_88_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_49_loopback_sample_req_88_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(41), ack => phi_stmt_49_req_1); -- 
    -- Element group access_T_CP_0_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_trigger
      -- 
    access_T_CP_0_elements(42) <= access_T_CP_0_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_entry_sample_req_ps
      -- 
    phi_stmt_49_entry_sample_req_91_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_49_entry_sample_req_91_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(43), ack => phi_stmt_49_req_0); -- 
    -- Element group access_T_CP_0_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_phi_mux_ack
      -- CP-element group 44: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_49_phi_mux_ack_ps
      -- 
    phi_stmt_49_phi_mux_ack_94_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_49_ack_0, ack => access_T_CP_0_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	49 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Sample/$entry
      -- CP-element group 47: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Sample/rr
      -- 
    rr_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(47), ack => type_cast_52_inst_req_0); -- 
    access_T_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(45) & access_T_CP_0_elements(49);
      gj_access_T_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_update_start_
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Update/cr
      -- 
    cr_112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(48), ack => type_cast_52_inst_req_1); -- 
    access_T_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(46) & access_T_CP_0_elements(50);
      gj_access_T_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	47 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Sample/ra
      -- 
    ra_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_0, ack => access_T_CP_0_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_update_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_52_Update/ca
      -- 
    ca_113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_52_inst_ack_1, ack => access_T_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_sample_start__ps
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Sample/req
      -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(51), ack => n_mycounter1_157_53_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_update_start__ps
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_update_start_
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Update/req
      -- 
    req_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(52), ack => n_mycounter1_157_53_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_sample_completed__ps
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Sample/ack
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter1_157_53_buf_ack_0, ack => access_T_CP_0_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_update_completed__ps
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter1_53_Update/ack
      -- 
    ack_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter1_157_53_buf_ack_1, ack => access_T_CP_0_elements(54)); -- 
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	12 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	11 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_start_
      -- 
    access_T_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	9 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	344 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	13 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_start_
      -- 
    access_T_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(344);
      gj_access_T_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	11 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_start__ps
      -- 
    access_T_CP_0_elements(57) <= access_T_CP_0_elements(11);
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	12 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	13 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_start__ps
      -- 
    access_T_CP_0_elements(59) <= access_T_CP_0_elements(13);
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	14 
    -- CP-element group 60: 	342 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	7 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_trigger
      -- 
    access_T_CP_0_elements(61) <= access_T_CP_0_elements(7);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_sample_req
      -- CP-element group 62: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_loopback_sample_req_ps
      -- 
    phi_stmt_54_loopback_sample_req_142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_54_loopback_sample_req_142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(62), ack => phi_stmt_54_req_1); -- 
    -- Element group access_T_CP_0_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	8 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_trigger
      -- 
    access_T_CP_0_elements(63) <= access_T_CP_0_elements(8);
    -- CP-element group 64:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_sample_req
      -- CP-element group 64: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_entry_sample_req_ps
      -- 
    phi_stmt_54_entry_sample_req_145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_54_entry_sample_req_145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(64), ack => phi_stmt_54_req_0); -- 
    -- Element group access_T_CP_0_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_phi_mux_ack
      -- CP-element group 65: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_54_phi_mux_ack_ps
      -- 
    phi_stmt_54_phi_mux_ack_148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_54_ack_0, ack => access_T_CP_0_elements(65)); -- 
    -- CP-element group 66:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_sample_start__ps
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_sample_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_update_start__ps
      -- CP-element group 67: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_update_start_
      -- 
    -- Element group access_T_CP_0_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_update_completed__ps
      -- 
    access_T_CP_0_elements(68) <= access_T_CP_0_elements(69);
    -- CP-element group 69:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	68 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_57_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(67), ack => access_T_CP_0_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Sample/req
      -- 
    req_169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(70), ack => n_row1_165_58_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_update_start__ps
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_update_start_
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Update/req
      -- 
    req_174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(71), ack => n_row1_165_58_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (4) 
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_sample_completed__ps
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Sample/ack
      -- 
    ack_170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_165_58_buf_ack_0, ack => access_T_CP_0_elements(72)); -- 
    -- CP-element group 73:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_update_completed__ps
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row1_58_Update/ack
      -- 
    ack_175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row1_165_58_buf_ack_1, ack => access_T_CP_0_elements(73)); -- 
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	9 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	12 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	11 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_start_
      -- 
    access_T_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	9 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	79 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	13 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_start_
      -- 
    access_T_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(79);
      gj_access_T_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	11 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_start__ps
      -- 
    access_T_CP_0_elements(76) <= access_T_CP_0_elements(11);
    -- CP-element group 77:  join  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	12 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	13 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_start__ps
      -- 
    access_T_CP_0_elements(78) <= access_T_CP_0_elements(13);
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	14 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	75 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	7 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_trigger
      -- 
    access_T_CP_0_elements(80) <= access_T_CP_0_elements(7);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_sample_req
      -- CP-element group 81: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_loopback_sample_req_ps
      -- 
    phi_stmt_59_loopback_sample_req_186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_loopback_sample_req_186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(81), ack => phi_stmt_59_req_0); -- 
    -- Element group access_T_CP_0_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	8 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_trigger
      -- 
    access_T_CP_0_elements(82) <= access_T_CP_0_elements(8);
    -- CP-element group 83:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_sample_req
      -- CP-element group 83: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_entry_sample_req_ps
      -- 
    phi_stmt_59_entry_sample_req_189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_59_entry_sample_req_189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(83), ack => phi_stmt_59_req_1); -- 
    -- Element group access_T_CP_0_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_phi_mux_ack
      -- CP-element group 84: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_59_phi_mux_ack_ps
      -- 
    phi_stmt_59_phi_mux_ack_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_59_ack_0, ack => access_T_CP_0_elements(84)); -- 
    -- CP-element group 85:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_sample_start__ps
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Sample/req
      -- 
    req_205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(85), ack => n_start1_146_61_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (4) 
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_update_start__ps
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_update_start_
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Update/req
      -- 
    req_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(86), ack => n_start1_146_61_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(86) is bound as output of CP function.
    -- CP-element group 87:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_sample_completed__ps
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_sample_completed_
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Sample/ack
      -- 
    ack_206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start1_146_61_buf_ack_0, ack => access_T_CP_0_elements(87)); -- 
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_update_completed__ps
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_update_completed_
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start1_61_Update/ack
      -- 
    ack_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start1_146_61_buf_ack_1, ack => access_T_CP_0_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_update_start__ps
      -- CP-element group 90: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_update_start_
      -- 
    -- Element group access_T_CP_0_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_update_completed__ps
      -- 
    access_T_CP_0_elements(91) <= access_T_CP_0_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_63_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(90), ack => access_T_CP_0_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  transition  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	9 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	12 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	11 
    -- CP-element group 93:  members (1) 
      -- CP-element group 93: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_sample_start_
      -- 
    access_T_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	9 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	352 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	13 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_update_start_
      -- 
    access_T_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "access_T_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(352);
      gj_access_T_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_sample_start__ps
      -- 
    access_T_CP_0_elements(95) <= access_T_CP_0_elements(11);
    -- CP-element group 96:  join  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	12 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(96) is bound as output of CP function.
    -- CP-element group 97:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	13 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_update_start__ps
      -- 
    access_T_CP_0_elements(97) <= access_T_CP_0_elements(13);
    -- CP-element group 98:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	14 
    -- CP-element group 98: 	352 
    -- CP-element group 98:  members (15) 
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_resize_1/index_resize_ack
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_resize_1/index_resize_req
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_resize_1/$exit
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_resize_1/$entry
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_computed_1
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_scaled_1
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_resized_1
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Sample/req
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_update_completed__ps
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_scale_1/scale_rename_ack
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_scale_1/scale_rename_req
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_scale_1/$exit
      -- CP-element group 98: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_index_scale_1/$entry
      -- 
    req_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(98), ack => array_obj_ref_203_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(98) is bound as output of CP function.
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	7 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_loopback_trigger
      -- 
    access_T_CP_0_elements(99) <= access_T_CP_0_elements(7);
    -- CP-element group 100:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_loopback_sample_req
      -- CP-element group 100: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_loopback_sample_req_ps
      -- 
    phi_stmt_64_loopback_sample_req_230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_64_loopback_sample_req_230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(100), ack => phi_stmt_64_req_0); -- 
    -- Element group access_T_CP_0_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	8 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_entry_trigger
      -- 
    access_T_CP_0_elements(101) <= access_T_CP_0_elements(8);
    -- CP-element group 102:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_entry_sample_req
      -- CP-element group 102: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_entry_sample_req_ps
      -- 
    phi_stmt_64_entry_sample_req_233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_64_entry_sample_req_233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(102), ack => phi_stmt_64_req_1); -- 
    -- Element group access_T_CP_0_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_phi_mux_ack
      -- CP-element group 103: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_64_phi_mux_ack_ps
      -- 
    phi_stmt_64_phi_mux_ack_236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_64_ack_0, ack => access_T_CP_0_elements(103)); -- 
    -- CP-element group 104:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_sample_start__ps
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_sample_start_
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Sample/$entry
      -- CP-element group 104: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Sample/req
      -- 
    req_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(104), ack => n_address2_241_66_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(104) is bound as output of CP function.
    -- CP-element group 105:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Update/$entry
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Update/req
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_update_start__ps
      -- CP-element group 105: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_update_start_
      -- 
    req_254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(105), ack => n_address2_241_66_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (4) 
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_sample_completed__ps
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Sample/ack
      -- 
    ack_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_241_66_buf_ack_0, ack => access_T_CP_0_elements(106)); -- 
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (4) 
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_Update/ack
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_update_completed__ps
      -- CP-element group 107: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address2_66_update_completed_
      -- 
    ack_255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_241_66_buf_ack_1, ack => access_T_CP_0_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: marked-predecessors 
    -- CP-element group 110: 	112 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_sample_start_
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Sample/$entry
      -- CP-element group 110: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Sample/rr
      -- 
    rr_267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(110), ack => type_cast_68_inst_req_0); -- 
    access_T_cp_element_group_110: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_110"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(108) & access_T_CP_0_elements(112);
      gj_access_T_cp_element_group_110 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(110), clk => clk, reset => reset); --
    end block;
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_update_start_
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Update/$entry
      -- CP-element group 111: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Update/cr
      -- 
    cr_272_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_272_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(111), ack => type_cast_68_inst_req_1); -- 
    access_T_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(109) & access_T_CP_0_elements(113);
      gj_access_T_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	110 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_sample_completed__ps
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Sample/ra
      -- 
    ra_268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_0, ack => access_T_CP_0_elements(112)); -- 
    -- CP-element group 113:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_update_completed__ps
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_68_Update/ca
      -- 
    ca_273_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_68_inst_ack_1, ack => access_T_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	9 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	12 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	11 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_sample_start_
      -- 
    access_T_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  join  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	9 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	119 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	13 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_update_start_
      -- 
    access_T_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(119);
      gj_access_T_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	11 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_sample_start__ps
      -- 
    access_T_CP_0_elements(116) <= access_T_CP_0_elements(11);
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	12 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(117) is bound as output of CP function.
    -- CP-element group 118:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	13 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_update_start__ps
      -- 
    access_T_CP_0_elements(118) <= access_T_CP_0_elements(13);
    -- CP-element group 119:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	14 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	115 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(119) is bound as output of CP function.
    -- CP-element group 120:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	7 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_loopback_trigger
      -- 
    access_T_CP_0_elements(120) <= access_T_CP_0_elements(7);
    -- CP-element group 121:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (2) 
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_loopback_sample_req
      -- CP-element group 121: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_loopback_sample_req_ps
      -- 
    phi_stmt_69_loopback_sample_req_284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_69_loopback_sample_req_284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(121), ack => phi_stmt_69_req_0); -- 
    -- Element group access_T_CP_0_elements(121) is bound as output of CP function.
    -- CP-element group 122:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	8 
    -- CP-element group 122: successors 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_entry_trigger
      -- 
    access_T_CP_0_elements(122) <= access_T_CP_0_elements(8);
    -- CP-element group 123:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: successors 
    -- CP-element group 123:  members (2) 
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_entry_sample_req
      -- CP-element group 123: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_entry_sample_req_ps
      -- 
    phi_stmt_69_entry_sample_req_287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_69_entry_sample_req_287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(123), ack => phi_stmt_69_req_1); -- 
    -- Element group access_T_CP_0_elements(123) is bound as output of CP function.
    -- CP-element group 124:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (2) 
      -- CP-element group 124: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_phi_mux_ack
      -- CP-element group 124: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_69_phi_mux_ack_ps
      -- 
    phi_stmt_69_phi_mux_ack_290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_69_ack_0, ack => access_T_CP_0_elements(124)); -- 
    -- CP-element group 125:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (4) 
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_sample_start__ps
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Sample/req
      -- 
    req_303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(125), ack => n_mycounter2_223_71_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(125) is bound as output of CP function.
    -- CP-element group 126:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (4) 
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_update_start__ps
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_update_start_
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Update/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(126), ack => n_mycounter2_223_71_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(126) is bound as output of CP function.
    -- CP-element group 127:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (4) 
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_sample_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Sample/ack
      -- 
    ack_304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter2_223_71_buf_ack_0, ack => access_T_CP_0_elements(127)); -- 
    -- CP-element group 128:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (4) 
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_update_completed__ps
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter2_71_Update/ack
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter2_223_71_buf_ack_1, ack => access_T_CP_0_elements(128)); -- 
    -- CP-element group 129:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	131 
    -- CP-element group 129:  members (1) 
      -- CP-element group 129: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(129) is bound as output of CP function.
    -- CP-element group 130:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(130) is bound as output of CP function.
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	129 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Sample/rr
      -- 
    rr_321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(131), ack => type_cast_73_inst_req_0); -- 
    access_T_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(129) & access_T_CP_0_elements(133);
      gj_access_T_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_update_start_
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Update/cr
      -- 
    cr_326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(132), ack => type_cast_73_inst_req_1); -- 
    access_T_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(130) & access_T_CP_0_elements(134);
      gj_access_T_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	131 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_sample_completed__ps
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Sample/ra
      -- 
    ra_322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_73_inst_ack_0, ack => access_T_CP_0_elements(133)); -- 
    -- CP-element group 134:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	132 
    -- CP-element group 134:  members (4) 
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_update_completed__ps
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_73_Update/ca
      -- 
    ca_327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_73_inst_ack_1, ack => access_T_CP_0_elements(134)); -- 
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	9 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	12 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	11 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_sample_start_
      -- 
    access_T_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	9 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	362 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	13 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_update_start_
      -- 
    access_T_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	11 
    -- CP-element group 137: successors 
    -- CP-element group 137:  members (1) 
      -- CP-element group 137: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_sample_start__ps
      -- 
    access_T_CP_0_elements(137) <= access_T_CP_0_elements(11);
    -- CP-element group 138:  join  transition  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	12 
    -- CP-element group 138:  members (1) 
      -- CP-element group 138: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(138) is bound as output of CP function.
    -- CP-element group 139:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	13 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (1) 
      -- CP-element group 139: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_update_start__ps
      -- 
    access_T_CP_0_elements(139) <= access_T_CP_0_elements(13);
    -- CP-element group 140:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	360 
    -- CP-element group 140: 	14 
    -- CP-element group 140:  members (2) 
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(140) is bound as output of CP function.
    -- CP-element group 141:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	7 
    -- CP-element group 141: successors 
    -- CP-element group 141:  members (1) 
      -- CP-element group 141: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_loopback_trigger
      -- 
    access_T_CP_0_elements(141) <= access_T_CP_0_elements(7);
    -- CP-element group 142:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: successors 
    -- CP-element group 142:  members (2) 
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_loopback_sample_req
      -- CP-element group 142: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_loopback_sample_req_ps
      -- 
    phi_stmt_74_loopback_sample_req_338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_loopback_sample_req_338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(142), ack => phi_stmt_74_req_1); -- 
    -- Element group access_T_CP_0_elements(142) is bound as output of CP function.
    -- CP-element group 143:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	8 
    -- CP-element group 143: successors 
    -- CP-element group 143:  members (1) 
      -- CP-element group 143: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_entry_trigger
      -- 
    access_T_CP_0_elements(143) <= access_T_CP_0_elements(8);
    -- CP-element group 144:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (2) 
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_entry_sample_req
      -- CP-element group 144: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_entry_sample_req_ps
      -- 
    phi_stmt_74_entry_sample_req_341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_74_entry_sample_req_341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(144), ack => phi_stmt_74_req_0); -- 
    -- Element group access_T_CP_0_elements(144) is bound as output of CP function.
    -- CP-element group 145:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: successors 
    -- CP-element group 145:  members (2) 
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_phi_mux_ack
      -- CP-element group 145: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_74_phi_mux_ack_ps
      -- 
    phi_stmt_74_phi_mux_ack_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_74_ack_0, ack => access_T_CP_0_elements(145)); -- 
    -- CP-element group 146:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: successors 
    -- CP-element group 146:  members (4) 
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_sample_start__ps
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_sample_completed__ps
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(146) is bound as output of CP function.
    -- CP-element group 147:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (2) 
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_update_start__ps
      -- CP-element group 147: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_update_start_
      -- 
    -- Element group access_T_CP_0_elements(147) is bound as output of CP function.
    -- CP-element group 148:  join  transition  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	149 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (1) 
      -- CP-element group 148: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_update_completed__ps
      -- 
    access_T_CP_0_elements(148) <= access_T_CP_0_elements(149);
    -- CP-element group 149:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	148 
    -- CP-element group 149:  members (1) 
      -- CP-element group 149: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_77_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(149) is a control-delay.
    cp_element_149_delay: control_delay_element  generic map(name => " 149_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(147), ack => access_T_CP_0_elements(149), clk => clk, reset =>reset);
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (4) 
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_sample_start__ps
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Sample/req
      -- 
    req_365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(150), ack => n_row2_231_78_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(150) is bound as output of CP function.
    -- CP-element group 151:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (4) 
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_update_start__ps
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_update_start_
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Update/req
      -- 
    req_370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(151), ack => n_row2_231_78_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(151) is bound as output of CP function.
    -- CP-element group 152:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (4) 
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_sample_completed__ps
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Sample/ack
      -- 
    ack_366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_231_78_buf_ack_0, ack => access_T_CP_0_elements(152)); -- 
    -- CP-element group 153:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153:  members (4) 
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_update_completed__ps
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row2_78_Update/ack
      -- 
    ack_371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row2_231_78_buf_ack_1, ack => access_T_CP_0_elements(153)); -- 
    -- CP-element group 154:  join  transition  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	9 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	12 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	11 
    -- CP-element group 154:  members (1) 
      -- CP-element group 154: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_sample_start_
      -- 
    access_T_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	9 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	159 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	13 
    -- CP-element group 155:  members (1) 
      -- CP-element group 155: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_update_start_
      -- 
    access_T_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(159);
      gj_access_T_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	11 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (1) 
      -- CP-element group 156: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_sample_start__ps
      -- 
    access_T_CP_0_elements(156) <= access_T_CP_0_elements(11);
    -- CP-element group 157:  join  transition  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	12 
    -- CP-element group 157:  members (1) 
      -- CP-element group 157: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(157) is bound as output of CP function.
    -- CP-element group 158:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	13 
    -- CP-element group 158: successors 
    -- CP-element group 158:  members (1) 
      -- CP-element group 158: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_update_start__ps
      -- 
    access_T_CP_0_elements(158) <= access_T_CP_0_elements(13);
    -- CP-element group 159:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	14 
    -- CP-element group 159: marked-successors 
    -- CP-element group 159: 	155 
    -- CP-element group 159:  members (2) 
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(159) is bound as output of CP function.
    -- CP-element group 160:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	7 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (1) 
      -- CP-element group 160: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_loopback_trigger
      -- 
    access_T_CP_0_elements(160) <= access_T_CP_0_elements(7);
    -- CP-element group 161:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: successors 
    -- CP-element group 161:  members (2) 
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_loopback_sample_req
      -- CP-element group 161: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_loopback_sample_req_ps
      -- 
    phi_stmt_79_loopback_sample_req_382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_79_loopback_sample_req_382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(161), ack => phi_stmt_79_req_1); -- 
    -- Element group access_T_CP_0_elements(161) is bound as output of CP function.
    -- CP-element group 162:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	8 
    -- CP-element group 162: successors 
    -- CP-element group 162:  members (1) 
      -- CP-element group 162: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_entry_trigger
      -- 
    access_T_CP_0_elements(162) <= access_T_CP_0_elements(8);
    -- CP-element group 163:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (2) 
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_entry_sample_req
      -- CP-element group 163: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_entry_sample_req_ps
      -- 
    phi_stmt_79_entry_sample_req_385_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_79_entry_sample_req_385_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(163), ack => phi_stmt_79_req_0); -- 
    -- Element group access_T_CP_0_elements(163) is bound as output of CP function.
    -- CP-element group 164:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (2) 
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_phi_mux_ack
      -- CP-element group 164: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_79_phi_mux_ack_ps
      -- 
    phi_stmt_79_phi_mux_ack_388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_79_ack_0, ack => access_T_CP_0_elements(164)); -- 
    -- CP-element group 165:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: successors 
    -- CP-element group 165:  members (4) 
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_sample_start__ps
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_sample_completed__ps
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(165) is bound as output of CP function.
    -- CP-element group 166:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (2) 
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_update_start__ps
      -- CP-element group 166: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_update_start_
      -- 
    -- Element group access_T_CP_0_elements(166) is bound as output of CP function.
    -- CP-element group 167:  join  transition  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	168 
    -- CP-element group 167: successors 
    -- CP-element group 167:  members (1) 
      -- CP-element group 167: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_update_completed__ps
      -- 
    access_T_CP_0_elements(167) <= access_T_CP_0_elements(168);
    -- CP-element group 168:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	167 
    -- CP-element group 168:  members (1) 
      -- CP-element group 168: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_82_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(168) is a control-delay.
    cp_element_168_delay: control_delay_element  generic map(name => " 168_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(166), ack => access_T_CP_0_elements(168), clk => clk, reset =>reset);
    -- CP-element group 169:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (4) 
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_sample_start__ps
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Sample/req
      -- 
    req_409_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_409_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(169), ack => n_start2_212_83_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(169) is bound as output of CP function.
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (4) 
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_update_start__ps
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_update_start_
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Update/req
      -- 
    req_414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(170), ack => n_start2_212_83_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(170) is bound as output of CP function.
    -- CP-element group 171:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (4) 
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_sample_completed__ps
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Sample/ack
      -- 
    ack_410_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start2_212_83_buf_ack_0, ack => access_T_CP_0_elements(171)); -- 
    -- CP-element group 172:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (4) 
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_update_completed__ps
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start2_83_Update/ack
      -- 
    ack_415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start2_212_83_buf_ack_1, ack => access_T_CP_0_elements(172)); -- 
    -- CP-element group 173:  join  transition  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	9 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	12 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	11 
    -- CP-element group 173:  members (1) 
      -- CP-element group 173: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_sample_start_
      -- 
    access_T_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	9 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	370 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	13 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_update_start_
      -- 
    access_T_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(370);
      gj_access_T_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	11 
    -- CP-element group 175: successors 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_sample_start__ps
      -- 
    access_T_CP_0_elements(175) <= access_T_CP_0_elements(11);
    -- CP-element group 176:  join  transition  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	12 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(176) is bound as output of CP function.
    -- CP-element group 177:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	13 
    -- CP-element group 177: successors 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_update_start__ps
      -- 
    access_T_CP_0_elements(177) <= access_T_CP_0_elements(13);
    -- CP-element group 178:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	370 
    -- CP-element group 178: 	14 
    -- CP-element group 178:  members (15) 
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/req
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_scale_1/scale_rename_ack
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_computed_1
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_resized_1
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_scale_1/scale_rename_req
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_resize_1/$entry
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_resize_1/$exit
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_scale_1/$entry
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_scale_1/$exit
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_scaled_1
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_resize_1/index_resize_ack
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_index_resize_1/index_resize_req
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_update_completed_
      -- CP-element group 178: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_update_completed__ps
      -- 
    req_1081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(178), ack => array_obj_ref_269_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(178) is bound as output of CP function.
    -- CP-element group 179:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	7 
    -- CP-element group 179: successors 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_loopback_trigger
      -- 
    access_T_CP_0_elements(179) <= access_T_CP_0_elements(7);
    -- CP-element group 180:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (2) 
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_loopback_sample_req
      -- CP-element group 180: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_loopback_sample_req_ps
      -- 
    phi_stmt_84_loopback_sample_req_426_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_84_loopback_sample_req_426_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(180), ack => phi_stmt_84_req_0); -- 
    -- Element group access_T_CP_0_elements(180) is bound as output of CP function.
    -- CP-element group 181:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	8 
    -- CP-element group 181: successors 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_entry_trigger
      -- 
    access_T_CP_0_elements(181) <= access_T_CP_0_elements(8);
    -- CP-element group 182:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_entry_sample_req
      -- CP-element group 182: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_entry_sample_req_ps
      -- 
    phi_stmt_84_entry_sample_req_429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_84_entry_sample_req_429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(182), ack => phi_stmt_84_req_1); -- 
    -- Element group access_T_CP_0_elements(182) is bound as output of CP function.
    -- CP-element group 183:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_phi_mux_ack
      -- CP-element group 183: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_84_phi_mux_ack_ps
      -- 
    phi_stmt_84_phi_mux_ack_432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_84_ack_0, ack => access_T_CP_0_elements(183)); -- 
    -- CP-element group 184:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (4) 
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_sample_start__ps
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_sample_start_
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Sample/$entry
      -- CP-element group 184: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Sample/req
      -- 
    req_445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(184), ack => n_address3_307_86_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(184) is bound as output of CP function.
    -- CP-element group 185:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (4) 
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_update_start__ps
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_update_start_
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Update/req
      -- 
    req_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(185), ack => n_address3_307_86_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(185) is bound as output of CP function.
    -- CP-element group 186:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (4) 
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_sample_completed__ps
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Sample/ack
      -- 
    ack_446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_307_86_buf_ack_0, ack => access_T_CP_0_elements(186)); -- 
    -- CP-element group 187:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187:  members (4) 
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_update_completed__ps
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address3_86_Update/ack
      -- 
    ack_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address3_307_86_buf_ack_1, ack => access_T_CP_0_elements(187)); -- 
    -- CP-element group 188:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (1) 
      -- CP-element group 188: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(188) is bound as output of CP function.
    -- CP-element group 189:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (1) 
      -- CP-element group 189: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(189) is bound as output of CP function.
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Sample/rr
      -- 
    rr_463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(190), ack => type_cast_88_inst_req_0); -- 
    access_T_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(188) & access_T_CP_0_elements(192);
      gj_access_T_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_update_start_
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Update/cr
      -- 
    cr_468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(191), ack => type_cast_88_inst_req_1); -- 
    access_T_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(189) & access_T_CP_0_elements(193);
      gj_access_T_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (4) 
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_sample_completed__ps
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Sample/ra
      -- 
    ra_464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_0, ack => access_T_CP_0_elements(192)); -- 
    -- CP-element group 193:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (4) 
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_update_completed__ps
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_88_Update/ca
      -- 
    ca_469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_88_inst_ack_1, ack => access_T_CP_0_elements(193)); -- 
    -- CP-element group 194:  join  transition  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	9 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	12 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	11 
    -- CP-element group 194:  members (1) 
      -- CP-element group 194: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_sample_start_
      -- 
    access_T_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	9 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	199 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	13 
    -- CP-element group 195:  members (1) 
      -- CP-element group 195: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_update_start_
      -- 
    access_T_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(199);
      gj_access_T_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	11 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (1) 
      -- CP-element group 196: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_sample_start__ps
      -- 
    access_T_CP_0_elements(196) <= access_T_CP_0_elements(11);
    -- CP-element group 197:  join  transition  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	12 
    -- CP-element group 197:  members (1) 
      -- CP-element group 197: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(197) is bound as output of CP function.
    -- CP-element group 198:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	13 
    -- CP-element group 198: successors 
    -- CP-element group 198:  members (1) 
      -- CP-element group 198: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_update_start__ps
      -- 
    access_T_CP_0_elements(198) <= access_T_CP_0_elements(13);
    -- CP-element group 199:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	14 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	195 
    -- CP-element group 199:  members (2) 
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(199) is bound as output of CP function.
    -- CP-element group 200:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	7 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (1) 
      -- CP-element group 200: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_loopback_trigger
      -- 
    access_T_CP_0_elements(200) <= access_T_CP_0_elements(7);
    -- CP-element group 201:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: successors 
    -- CP-element group 201:  members (2) 
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_loopback_sample_req
      -- CP-element group 201: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_loopback_sample_req_ps
      -- 
    phi_stmt_89_loopback_sample_req_480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_89_loopback_sample_req_480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(201), ack => phi_stmt_89_req_0); -- 
    -- Element group access_T_CP_0_elements(201) is bound as output of CP function.
    -- CP-element group 202:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	8 
    -- CP-element group 202: successors 
    -- CP-element group 202:  members (1) 
      -- CP-element group 202: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_entry_trigger
      -- 
    access_T_CP_0_elements(202) <= access_T_CP_0_elements(8);
    -- CP-element group 203:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: successors 
    -- CP-element group 203:  members (2) 
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_entry_sample_req
      -- CP-element group 203: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_entry_sample_req_ps
      -- 
    phi_stmt_89_entry_sample_req_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_89_entry_sample_req_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(203), ack => phi_stmt_89_req_1); -- 
    -- Element group access_T_CP_0_elements(203) is bound as output of CP function.
    -- CP-element group 204:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (2) 
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_phi_mux_ack
      -- CP-element group 204: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_89_phi_mux_ack_ps
      -- 
    phi_stmt_89_phi_mux_ack_486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_89_ack_0, ack => access_T_CP_0_elements(204)); -- 
    -- CP-element group 205:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	207 
    -- CP-element group 205:  members (4) 
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_sample_start__ps
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Sample/req
      -- 
    req_499_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_499_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(205), ack => n_mycounter3_289_91_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(205) is bound as output of CP function.
    -- CP-element group 206:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (4) 
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_update_start__ps
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_update_start_
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Update/req
      -- 
    req_504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(206), ack => n_mycounter3_289_91_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(206) is bound as output of CP function.
    -- CP-element group 207:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	205 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (4) 
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_sample_completed__ps
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Sample/$exit
      -- CP-element group 207: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Sample/ack
      -- 
    ack_500_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter3_289_91_buf_ack_0, ack => access_T_CP_0_elements(207)); -- 
    -- CP-element group 208:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208:  members (4) 
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_update_completed__ps
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_update_completed_
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter3_91_Update/ack
      -- 
    ack_505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter3_289_91_buf_ack_1, ack => access_T_CP_0_elements(208)); -- 
    -- CP-element group 209:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (1) 
      -- CP-element group 209: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(209) is bound as output of CP function.
    -- CP-element group 210:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (1) 
      -- CP-element group 210: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(210) is bound as output of CP function.
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_sample_start_
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Sample/rr
      -- 
    rr_517_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_517_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(211), ack => type_cast_93_inst_req_0); -- 
    access_T_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(209) & access_T_CP_0_elements(213);
      gj_access_T_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: marked-predecessors 
    -- CP-element group 212: 	214 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	214 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_update_start_
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Update/$entry
      -- CP-element group 212: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Update/cr
      -- 
    cr_522_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_522_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(212), ack => type_cast_93_inst_req_1); -- 
    access_T_cp_element_group_212: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_212"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(210) & access_T_CP_0_elements(214);
      gj_access_T_cp_element_group_212 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(212), clk => clk, reset => reset); --
    end block;
    -- CP-element group 213:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (4) 
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_sample_completed__ps
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_sample_completed_
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Sample/$exit
      -- CP-element group 213: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Sample/ra
      -- 
    ra_518_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_0, ack => access_T_CP_0_elements(213)); -- 
    -- CP-element group 214:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	212 
    -- CP-element group 214: successors 
    -- CP-element group 214: marked-successors 
    -- CP-element group 214: 	212 
    -- CP-element group 214:  members (4) 
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_update_completed__ps
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_update_completed_
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Update/$exit
      -- CP-element group 214: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_93_Update/ca
      -- 
    ca_523_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_93_inst_ack_1, ack => access_T_CP_0_elements(214)); -- 
    -- CP-element group 215:  join  transition  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	9 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	12 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	11 
    -- CP-element group 215:  members (1) 
      -- CP-element group 215: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_sample_start_
      -- 
    access_T_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  join  transition  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	9 
    -- CP-element group 216: marked-predecessors 
    -- CP-element group 216: 	380 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	13 
    -- CP-element group 216:  members (1) 
      -- CP-element group 216: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_update_start_
      -- 
    access_T_cp_element_group_216: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_216"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(380);
      gj_access_T_cp_element_group_216 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(216), clk => clk, reset => reset); --
    end block;
    -- CP-element group 217:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	11 
    -- CP-element group 217: successors 
    -- CP-element group 217:  members (1) 
      -- CP-element group 217: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_sample_start__ps
      -- 
    access_T_CP_0_elements(217) <= access_T_CP_0_elements(11);
    -- CP-element group 218:  join  transition  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	12 
    -- CP-element group 218:  members (1) 
      -- CP-element group 218: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(218) is bound as output of CP function.
    -- CP-element group 219:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	13 
    -- CP-element group 219: successors 
    -- CP-element group 219:  members (1) 
      -- CP-element group 219: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_update_start__ps
      -- 
    access_T_CP_0_elements(219) <= access_T_CP_0_elements(13);
    -- CP-element group 220:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	378 
    -- CP-element group 220: 	14 
    -- CP-element group 220:  members (2) 
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(220) is bound as output of CP function.
    -- CP-element group 221:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	7 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (1) 
      -- CP-element group 221: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_loopback_trigger
      -- 
    access_T_CP_0_elements(221) <= access_T_CP_0_elements(7);
    -- CP-element group 222:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: successors 
    -- CP-element group 222:  members (2) 
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_loopback_sample_req
      -- CP-element group 222: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_loopback_sample_req_ps
      -- 
    phi_stmt_94_loopback_sample_req_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_94_loopback_sample_req_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(222), ack => phi_stmt_94_req_1); -- 
    -- Element group access_T_CP_0_elements(222) is bound as output of CP function.
    -- CP-element group 223:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	8 
    -- CP-element group 223: successors 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_entry_trigger
      -- 
    access_T_CP_0_elements(223) <= access_T_CP_0_elements(8);
    -- CP-element group 224:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_entry_sample_req
      -- CP-element group 224: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_entry_sample_req_ps
      -- 
    phi_stmt_94_entry_sample_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_94_entry_sample_req_537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(224), ack => phi_stmt_94_req_0); -- 
    -- Element group access_T_CP_0_elements(224) is bound as output of CP function.
    -- CP-element group 225:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_phi_mux_ack
      -- CP-element group 225: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_94_phi_mux_ack_ps
      -- 
    phi_stmt_94_phi_mux_ack_540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_94_ack_0, ack => access_T_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: successors 
    -- CP-element group 226:  members (4) 
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_sample_start__ps
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_sample_completed__ps
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(226) is bound as output of CP function.
    -- CP-element group 227:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (2) 
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_update_start__ps
      -- CP-element group 227: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_update_start_
      -- 
    -- Element group access_T_CP_0_elements(227) is bound as output of CP function.
    -- CP-element group 228:  join  transition  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	229 
    -- CP-element group 228: successors 
    -- CP-element group 228:  members (1) 
      -- CP-element group 228: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_update_completed__ps
      -- 
    access_T_CP_0_elements(228) <= access_T_CP_0_elements(229);
    -- CP-element group 229:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	228 
    -- CP-element group 229:  members (1) 
      -- CP-element group 229: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_97_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(229) is a control-delay.
    cp_element_229_delay: control_delay_element  generic map(name => " 229_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(227), ack => access_T_CP_0_elements(229), clk => clk, reset =>reset);
    -- CP-element group 230:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (4) 
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_sample_start__ps
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Sample/req
      -- 
    req_561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(230), ack => n_row3_297_98_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(230) is bound as output of CP function.
    -- CP-element group 231:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (4) 
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_update_start__ps
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_update_start_
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Update/req
      -- 
    req_566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(231), ack => n_row3_297_98_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(231) is bound as output of CP function.
    -- CP-element group 232:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (4) 
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_sample_completed__ps
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Sample/ack
      -- 
    ack_562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_297_98_buf_ack_0, ack => access_T_CP_0_elements(232)); -- 
    -- CP-element group 233:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (4) 
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_update_completed__ps
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row3_98_Update/ack
      -- 
    ack_567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row3_297_98_buf_ack_1, ack => access_T_CP_0_elements(233)); -- 
    -- CP-element group 234:  join  transition  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	9 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	12 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	11 
    -- CP-element group 234:  members (1) 
      -- CP-element group 234: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_sample_start_
      -- 
    access_T_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	9 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	239 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	13 
    -- CP-element group 235:  members (1) 
      -- CP-element group 235: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_update_start_
      -- 
    access_T_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(239);
      gj_access_T_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	11 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (1) 
      -- CP-element group 236: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_sample_start__ps
      -- 
    access_T_CP_0_elements(236) <= access_T_CP_0_elements(11);
    -- CP-element group 237:  join  transition  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	12 
    -- CP-element group 237:  members (1) 
      -- CP-element group 237: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(237) is bound as output of CP function.
    -- CP-element group 238:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	13 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (1) 
      -- CP-element group 238: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_update_start__ps
      -- 
    access_T_CP_0_elements(238) <= access_T_CP_0_elements(13);
    -- CP-element group 239:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	14 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	235 
    -- CP-element group 239:  members (2) 
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(239) is bound as output of CP function.
    -- CP-element group 240:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	7 
    -- CP-element group 240: successors 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_loopback_trigger
      -- 
    access_T_CP_0_elements(240) <= access_T_CP_0_elements(7);
    -- CP-element group 241:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (2) 
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_loopback_sample_req
      -- CP-element group 241: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_loopback_sample_req_ps
      -- 
    phi_stmt_99_loopback_sample_req_578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_99_loopback_sample_req_578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(241), ack => phi_stmt_99_req_0); -- 
    -- Element group access_T_CP_0_elements(241) is bound as output of CP function.
    -- CP-element group 242:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	8 
    -- CP-element group 242: successors 
    -- CP-element group 242:  members (1) 
      -- CP-element group 242: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_entry_trigger
      -- 
    access_T_CP_0_elements(242) <= access_T_CP_0_elements(8);
    -- CP-element group 243:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: successors 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_entry_sample_req
      -- CP-element group 243: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_entry_sample_req_ps
      -- 
    phi_stmt_99_entry_sample_req_581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_99_entry_sample_req_581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(243), ack => phi_stmt_99_req_1); -- 
    -- Element group access_T_CP_0_elements(243) is bound as output of CP function.
    -- CP-element group 244:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (2) 
      -- CP-element group 244: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_phi_mux_ack
      -- CP-element group 244: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_99_phi_mux_ack_ps
      -- 
    phi_stmt_99_phi_mux_ack_584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_99_ack_0, ack => access_T_CP_0_elements(244)); -- 
    -- CP-element group 245:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (4) 
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_sample_start__ps
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Sample/req
      -- 
    req_597_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_597_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(245), ack => n_start3_278_101_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(245) is bound as output of CP function.
    -- CP-element group 246:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (4) 
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_update_start__ps
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_update_start_
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Update/req
      -- 
    req_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(246), ack => n_start3_278_101_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(246) is bound as output of CP function.
    -- CP-element group 247:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247:  members (4) 
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_sample_completed__ps
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Sample/ack
      -- 
    ack_598_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start3_278_101_buf_ack_0, ack => access_T_CP_0_elements(247)); -- 
    -- CP-element group 248:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (4) 
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_update_completed__ps
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start3_101_Update/ack
      -- 
    ack_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start3_278_101_buf_ack_1, ack => access_T_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: successors 
    -- CP-element group 249:  members (4) 
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_sample_start__ps
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_sample_completed__ps
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_sample_completed_
      -- 
    -- Element group access_T_CP_0_elements(249) is bound as output of CP function.
    -- CP-element group 250:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_update_start__ps
      -- CP-element group 250: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_update_start_
      -- 
    -- Element group access_T_CP_0_elements(250) is bound as output of CP function.
    -- CP-element group 251:  join  transition  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	252 
    -- CP-element group 251: successors 
    -- CP-element group 251:  members (1) 
      -- CP-element group 251: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_update_completed__ps
      -- 
    access_T_CP_0_elements(251) <= access_T_CP_0_elements(252);
    -- CP-element group 252:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	251 
    -- CP-element group 252:  members (1) 
      -- CP-element group 252: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_103_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(252) is a control-delay.
    cp_element_252_delay: control_delay_element  generic map(name => " 252_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(250), ack => access_T_CP_0_elements(252), clk => clk, reset =>reset);
    -- CP-element group 253:  join  transition  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	9 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	12 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	11 
    -- CP-element group 253:  members (1) 
      -- CP-element group 253: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_sample_start_
      -- 
    access_T_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	9 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	388 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	13 
    -- CP-element group 254:  members (1) 
      -- CP-element group 254: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_update_start_
      -- 
    access_T_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(388);
      gj_access_T_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	11 
    -- CP-element group 255: successors 
    -- CP-element group 255:  members (1) 
      -- CP-element group 255: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_sample_start__ps
      -- 
    access_T_CP_0_elements(255) <= access_T_CP_0_elements(11);
    -- CP-element group 256:  join  transition  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	12 
    -- CP-element group 256:  members (1) 
      -- CP-element group 256: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(256) is bound as output of CP function.
    -- CP-element group 257:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	13 
    -- CP-element group 257: successors 
    -- CP-element group 257:  members (1) 
      -- CP-element group 257: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_update_start__ps
      -- 
    access_T_CP_0_elements(257) <= access_T_CP_0_elements(13);
    -- CP-element group 258:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	388 
    -- CP-element group 258: 	14 
    -- CP-element group 258:  members (15) 
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_update_completed_
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_update_completed__ps
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_resized_1
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_scaled_1
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_computed_1
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_resize_1/$entry
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_resize_1/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_resize_1/index_resize_req
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_resize_1/index_resize_ack
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_scale_1/$entry
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_scale_1/$exit
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_scale_1/scale_rename_req
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_index_scale_1/scale_rename_ack
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Sample/req
      -- 
    req_1205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(258), ack => array_obj_ref_335_index_offset_req_0); -- 
    -- Element group access_T_CP_0_elements(258) is bound as output of CP function.
    -- CP-element group 259:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	7 
    -- CP-element group 259: successors 
    -- CP-element group 259:  members (1) 
      -- CP-element group 259: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_loopback_trigger
      -- 
    access_T_CP_0_elements(259) <= access_T_CP_0_elements(7);
    -- CP-element group 260:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: successors 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_loopback_sample_req
      -- CP-element group 260: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_loopback_sample_req_ps
      -- 
    phi_stmt_104_loopback_sample_req_622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_104_loopback_sample_req_622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(260), ack => phi_stmt_104_req_1); -- 
    -- Element group access_T_CP_0_elements(260) is bound as output of CP function.
    -- CP-element group 261:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	8 
    -- CP-element group 261: successors 
    -- CP-element group 261:  members (1) 
      -- CP-element group 261: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_entry_trigger
      -- 
    access_T_CP_0_elements(261) <= access_T_CP_0_elements(8);
    -- CP-element group 262:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: successors 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_entry_sample_req
      -- CP-element group 262: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_entry_sample_req_ps
      -- 
    phi_stmt_104_entry_sample_req_625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_104_entry_sample_req_625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(262), ack => phi_stmt_104_req_0); -- 
    -- Element group access_T_CP_0_elements(262) is bound as output of CP function.
    -- CP-element group 263:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: successors 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_phi_mux_ack
      -- CP-element group 263: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_104_phi_mux_ack_ps
      -- 
    phi_stmt_104_phi_mux_ack_628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_104_ack_0, ack => access_T_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (1) 
      -- CP-element group 264: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(264) is bound as output of CP function.
    -- CP-element group 265:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (1) 
      -- CP-element group 265: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(265) is bound as output of CP function.
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Sample/rr
      -- 
    rr_641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(266), ack => type_cast_109_inst_req_0); -- 
    access_T_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(264) & access_T_CP_0_elements(268);
      gj_access_T_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	269 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_start_
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Update/cr
      -- 
    cr_646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(267), ack => type_cast_109_inst_req_1); -- 
    access_T_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(265) & access_T_CP_0_elements(269);
      gj_access_T_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (4) 
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_completed__ps
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Sample/ra
      -- 
    ra_642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_109_inst_ack_0, ack => access_T_CP_0_elements(268)); -- 
    -- CP-element group 269:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: marked-successors 
    -- CP-element group 269: 	267 
    -- CP-element group 269:  members (4) 
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_completed__ps
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_109_Update/ca
      -- 
    ca_647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_109_inst_ack_1, ack => access_T_CP_0_elements(269)); -- 
    -- CP-element group 270:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (4) 
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_sample_start__ps
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Sample/req
      -- 
    req_659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(270), ack => n_address4_373_110_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(270) is bound as output of CP function.
    -- CP-element group 271:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (4) 
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_update_start__ps
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_update_start_
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Update/req
      -- 
    req_664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(271), ack => n_address4_373_110_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(271) is bound as output of CP function.
    -- CP-element group 272:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272:  members (4) 
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_sample_completed__ps
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Sample/ack
      -- 
    ack_660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_373_110_buf_ack_0, ack => access_T_CP_0_elements(272)); -- 
    -- CP-element group 273:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273:  members (4) 
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_update_completed__ps
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_address4_110_Update/ack
      -- 
    ack_665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address4_373_110_buf_ack_1, ack => access_T_CP_0_elements(273)); -- 
    -- CP-element group 274:  join  transition  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	9 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	12 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	11 
    -- CP-element group 274:  members (1) 
      -- CP-element group 274: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_start_
      -- 
    access_T_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  join  transition  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	9 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	279 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	13 
    -- CP-element group 275:  members (1) 
      -- CP-element group 275: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_start_
      -- 
    access_T_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(279);
      gj_access_T_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	11 
    -- CP-element group 276: successors 
    -- CP-element group 276:  members (1) 
      -- CP-element group 276: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_start__ps
      -- 
    access_T_CP_0_elements(276) <= access_T_CP_0_elements(11);
    -- CP-element group 277:  join  transition  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	12 
    -- CP-element group 277:  members (1) 
      -- CP-element group 277: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(277) is bound as output of CP function.
    -- CP-element group 278:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	13 
    -- CP-element group 278: successors 
    -- CP-element group 278:  members (1) 
      -- CP-element group 278: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_start__ps
      -- 
    access_T_CP_0_elements(278) <= access_T_CP_0_elements(13);
    -- CP-element group 279:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	14 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	275 
    -- CP-element group 279:  members (2) 
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(279) is bound as output of CP function.
    -- CP-element group 280:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	7 
    -- CP-element group 280: successors 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_trigger
      -- 
    access_T_CP_0_elements(280) <= access_T_CP_0_elements(7);
    -- CP-element group 281:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: successors 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_sample_req
      -- CP-element group 281: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_loopback_sample_req_ps
      -- 
    phi_stmt_111_loopback_sample_req_676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_loopback_sample_req_676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(281), ack => phi_stmt_111_req_0); -- 
    -- Element group access_T_CP_0_elements(281) is bound as output of CP function.
    -- CP-element group 282:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	8 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_trigger
      -- 
    access_T_CP_0_elements(282) <= access_T_CP_0_elements(8);
    -- CP-element group 283:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: successors 
    -- CP-element group 283:  members (2) 
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_sample_req
      -- CP-element group 283: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_entry_sample_req_ps
      -- 
    phi_stmt_111_entry_sample_req_679_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_111_entry_sample_req_679_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(283), ack => phi_stmt_111_req_1); -- 
    -- Element group access_T_CP_0_elements(283) is bound as output of CP function.
    -- CP-element group 284:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: successors 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_phi_mux_ack
      -- CP-element group 284: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_111_phi_mux_ack_ps
      -- 
    phi_stmt_111_phi_mux_ack_682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_111_ack_0, ack => access_T_CP_0_elements(284)); -- 
    -- CP-element group 285:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (4) 
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_sample_start__ps
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Sample/req
      -- 
    req_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(285), ack => n_mycounter4_355_113_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(285) is bound as output of CP function.
    -- CP-element group 286:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (4) 
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_update_start__ps
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_update_start_
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Update/req
      -- 
    req_700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(286), ack => n_mycounter4_355_113_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(286) is bound as output of CP function.
    -- CP-element group 287:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287:  members (4) 
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_sample_completed__ps
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Sample/ack
      -- 
    ack_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter4_355_113_buf_ack_0, ack => access_T_CP_0_elements(287)); -- 
    -- CP-element group 288:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288:  members (4) 
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_update_completed__ps
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Update/$exit
      -- CP-element group 288: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_mycounter4_113_Update/ack
      -- 
    ack_701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_mycounter4_355_113_buf_ack_1, ack => access_T_CP_0_elements(288)); -- 
    -- CP-element group 289:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (1) 
      -- CP-element group 289: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(289) is bound as output of CP function.
    -- CP-element group 290:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (1) 
      -- CP-element group 290: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(290) is bound as output of CP function.
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	293 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_sample_start_
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Sample/$entry
      -- CP-element group 291: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Sample/rr
      -- 
    rr_713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(291), ack => type_cast_115_inst_req_0); -- 
    access_T_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(289) & access_T_CP_0_elements(293);
      gj_access_T_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: marked-predecessors 
    -- CP-element group 292: 	294 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	294 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_update_start_
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Update/$entry
      -- CP-element group 292: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Update/cr
      -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(292), ack => type_cast_115_inst_req_1); -- 
    access_T_cp_element_group_292: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_292"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(290) & access_T_CP_0_elements(294);
      gj_access_T_cp_element_group_292 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(292), clk => clk, reset => reset); --
    end block;
    -- CP-element group 293:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: marked-successors 
    -- CP-element group 293: 	291 
    -- CP-element group 293:  members (4) 
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_sample_completed__ps
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_sample_completed_
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Sample/$exit
      -- CP-element group 293: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Sample/ra
      -- 
    ra_714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_0, ack => access_T_CP_0_elements(293)); -- 
    -- CP-element group 294:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	292 
    -- CP-element group 294: successors 
    -- CP-element group 294: marked-successors 
    -- CP-element group 294: 	292 
    -- CP-element group 294:  members (4) 
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_update_completed__ps
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_update_completed_
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Update/$exit
      -- CP-element group 294: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_115_Update/ca
      -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 294_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_115_inst_ack_1, ack => access_T_CP_0_elements(294)); -- 
    -- CP-element group 295:  join  transition  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	9 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	12 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	11 
    -- CP-element group 295:  members (1) 
      -- CP-element group 295: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_start_
      -- 
    access_T_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  join  transition  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	9 
    -- CP-element group 296: marked-predecessors 
    -- CP-element group 296: 	398 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	13 
    -- CP-element group 296:  members (1) 
      -- CP-element group 296: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_start_
      -- 
    access_T_cp_element_group_296: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_296"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(398);
      gj_access_T_cp_element_group_296 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(296), clk => clk, reset => reset); --
    end block;
    -- CP-element group 297:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	11 
    -- CP-element group 297: successors 
    -- CP-element group 297:  members (1) 
      -- CP-element group 297: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_start__ps
      -- 
    access_T_CP_0_elements(297) <= access_T_CP_0_elements(11);
    -- CP-element group 298:  join  transition  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	12 
    -- CP-element group 298:  members (1) 
      -- CP-element group 298: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(298) is bound as output of CP function.
    -- CP-element group 299:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	13 
    -- CP-element group 299: successors 
    -- CP-element group 299:  members (1) 
      -- CP-element group 299: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_start__ps
      -- 
    access_T_CP_0_elements(299) <= access_T_CP_0_elements(13);
    -- CP-element group 300:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	396 
    -- CP-element group 300: 	14 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(300) is bound as output of CP function.
    -- CP-element group 301:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	7 
    -- CP-element group 301: successors 
    -- CP-element group 301:  members (1) 
      -- CP-element group 301: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_trigger
      -- 
    access_T_CP_0_elements(301) <= access_T_CP_0_elements(7);
    -- CP-element group 302:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: successors 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_sample_req_ps
      -- CP-element group 302: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_loopback_sample_req
      -- 
    phi_stmt_116_loopback_sample_req_730_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_loopback_sample_req_730_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(302), ack => phi_stmt_116_req_1); -- 
    -- Element group access_T_CP_0_elements(302) is bound as output of CP function.
    -- CP-element group 303:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	8 
    -- CP-element group 303: successors 
    -- CP-element group 303:  members (1) 
      -- CP-element group 303: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_trigger
      -- 
    access_T_CP_0_elements(303) <= access_T_CP_0_elements(8);
    -- CP-element group 304:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: successors 
    -- CP-element group 304:  members (2) 
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_sample_req_ps
      -- CP-element group 304: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_entry_sample_req
      -- 
    phi_stmt_116_entry_sample_req_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_116_entry_sample_req_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(304), ack => phi_stmt_116_req_0); -- 
    -- Element group access_T_CP_0_elements(304) is bound as output of CP function.
    -- CP-element group 305:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: successors 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_phi_mux_ack_ps
      -- CP-element group 305: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_116_phi_mux_ack
      -- 
    phi_stmt_116_phi_mux_ack_736_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_116_ack_0, ack => access_T_CP_0_elements(305)); -- 
    -- CP-element group 306:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: successors 
    -- CP-element group 306:  members (4) 
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_completed_
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_completed__ps
      -- CP-element group 306: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(306) is bound as output of CP function.
    -- CP-element group 307:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (2) 
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_start_
      -- CP-element group 307: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(307) is bound as output of CP function.
    -- CP-element group 308:  join  transition  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	309 
    -- CP-element group 308: successors 
    -- CP-element group 308:  members (1) 
      -- CP-element group 308: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_completed__ps
      -- 
    access_T_CP_0_elements(308) <= access_T_CP_0_elements(309);
    -- CP-element group 309:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	308 
    -- CP-element group 309:  members (1) 
      -- CP-element group 309: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_119_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(309) is a control-delay.
    cp_element_309_delay: control_delay_element  generic map(name => " 309_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(307), ack => access_T_CP_0_elements(309), clk => clk, reset =>reset);
    -- CP-element group 310:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (4) 
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_sample_start__ps
      -- 
    req_757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(310), ack => n_row4_363_120_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(310) is bound as output of CP function.
    -- CP-element group 311:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (4) 
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Update/req
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_update_start_
      -- CP-element group 311: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_update_start__ps
      -- 
    req_762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(311), ack => n_row4_363_120_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(311) is bound as output of CP function.
    -- CP-element group 312:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312:  members (4) 
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_sample_completed_
      -- CP-element group 312: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_sample_completed__ps
      -- 
    ack_758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row4_363_120_buf_ack_0, ack => access_T_CP_0_elements(312)); -- 
    -- CP-element group 313:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313:  members (4) 
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_update_completed_
      -- CP-element group 313: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_row4_120_update_completed__ps
      -- 
    ack_763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row4_363_120_buf_ack_1, ack => access_T_CP_0_elements(313)); -- 
    -- CP-element group 314:  join  transition  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	9 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	12 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	11 
    -- CP-element group 314:  members (1) 
      -- CP-element group 314: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_start_
      -- 
    access_T_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(12);
      gj_access_T_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  join  transition  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	9 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	317 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	13 
    -- CP-element group 315:  members (1) 
      -- CP-element group 315: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_start_
      -- 
    access_T_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(317);
      gj_access_T_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  join  transition  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	12 
    -- CP-element group 316:  members (1) 
      -- CP-element group 316: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_sample_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(316) is bound as output of CP function.
    -- CP-element group 317:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	14 
    -- CP-element group 317: marked-successors 
    -- CP-element group 317: 	315 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_completed_
      -- CP-element group 317: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_update_completed__ps
      -- 
    -- Element group access_T_CP_0_elements(317) is bound as output of CP function.
    -- CP-element group 318:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	7 
    -- CP-element group 318: successors 
    -- CP-element group 318:  members (1) 
      -- CP-element group 318: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_trigger
      -- 
    access_T_CP_0_elements(318) <= access_T_CP_0_elements(7);
    -- CP-element group 319:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: successors 
    -- CP-element group 319:  members (2) 
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_sample_req_ps
      -- CP-element group 319: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_loopback_sample_req
      -- 
    phi_stmt_121_loopback_sample_req_774_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_121_loopback_sample_req_774_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(319), ack => phi_stmt_121_req_0); -- 
    -- Element group access_T_CP_0_elements(319) is bound as output of CP function.
    -- CP-element group 320:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	8 
    -- CP-element group 320: successors 
    -- CP-element group 320:  members (1) 
      -- CP-element group 320: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_trigger
      -- 
    access_T_CP_0_elements(320) <= access_T_CP_0_elements(8);
    -- CP-element group 321:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: successors 
    -- CP-element group 321:  members (2) 
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_sample_req_ps
      -- CP-element group 321: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_entry_sample_req
      -- 
    phi_stmt_121_entry_sample_req_777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_121_entry_sample_req_777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(321), ack => phi_stmt_121_req_1); -- 
    -- Element group access_T_CP_0_elements(321) is bound as output of CP function.
    -- CP-element group 322:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: successors 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_phi_mux_ack_ps
      -- CP-element group 322: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/phi_stmt_121_phi_mux_ack
      -- 
    phi_stmt_121_phi_mux_ack_780_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_121_ack_0, ack => access_T_CP_0_elements(322)); -- 
    -- CP-element group 323:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (4) 
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Sample/req
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Sample/$entry
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_sample_start_
      -- CP-element group 323: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_sample_start__ps
      -- 
    req_793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(323), ack => n_start4_344_123_buf_req_0); -- 
    -- Element group access_T_CP_0_elements(323) is bound as output of CP function.
    -- CP-element group 324:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	326 
    -- CP-element group 324:  members (4) 
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Update/req
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Update/$entry
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_update_start_
      -- CP-element group 324: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_update_start__ps
      -- 
    req_798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(324), ack => n_start4_344_123_buf_req_1); -- 
    -- Element group access_T_CP_0_elements(324) is bound as output of CP function.
    -- CP-element group 325:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325:  members (4) 
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Sample/ack
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Sample/$exit
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_sample_completed_
      -- CP-element group 325: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_sample_completed__ps
      -- 
    ack_794_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start4_344_123_buf_ack_0, ack => access_T_CP_0_elements(325)); -- 
    -- CP-element group 326:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	324 
    -- CP-element group 326: successors 
    -- CP-element group 326:  members (4) 
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Update/$exit
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_update_completed_
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_update_completed__ps
      -- CP-element group 326: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/R_n_start4_123_Update/ack
      -- 
    ack_799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_start4_344_123_buf_ack_1, ack => access_T_CP_0_elements(326)); -- 
    -- CP-element group 327:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: successors 
    -- CP-element group 327:  members (4) 
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_sample_start_
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_sample_completed__ps
      -- CP-element group 327: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_sample_start__ps
      -- 
    -- Element group access_T_CP_0_elements(327) is bound as output of CP function.
    -- CP-element group 328:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	330 
    -- CP-element group 328:  members (2) 
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_update_start_
      -- CP-element group 328: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_update_start__ps
      -- 
    -- Element group access_T_CP_0_elements(328) is bound as output of CP function.
    -- CP-element group 329:  join  transition  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	330 
    -- CP-element group 329: successors 
    -- CP-element group 329:  members (1) 
      -- CP-element group 329: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_update_completed__ps
      -- 
    access_T_CP_0_elements(329) <= access_T_CP_0_elements(330);
    -- CP-element group 330:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	328 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	329 
    -- CP-element group 330:  members (1) 
      -- CP-element group 330: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/type_cast_125_update_completed_
      -- 
    -- Element group access_T_CP_0_elements(330) is a control-delay.
    cp_element_330_delay: control_delay_element  generic map(name => " 330_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(328), ack => access_T_CP_0_elements(330), clk => clk, reset =>reset);
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	335 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	336 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	336 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_request/req
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_request/$entry
      -- CP-element group 331: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_sample_start_
      -- 
    req_848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(331), ack => addr_of_138_final_reg_req_0); -- 
    access_T_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(335) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	9 
    -- CP-element group 332: marked-predecessors 
    -- CP-element group 332: 	340 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	337 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_complete/req
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_complete/$entry
      -- CP-element group 332: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_update_start_
      -- 
    req_853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(332), ack => addr_of_138_final_reg_req_1); -- 
    access_T_cp_element_group_332: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_332"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(340);
      gj_access_T_cp_element_group_332 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(332), clk => clk, reset => reset); --
    end block;
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	9 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	336 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Update/req
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Update/$entry
      -- CP-element group 333: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_update_start
      -- 
    req_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(333), ack => array_obj_ref_137_index_offset_req_1); -- 
    access_T_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(336);
      gj_access_T_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	20 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	404 
    -- CP-element group 334: marked-successors 
    -- CP-element group 334: 	16 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Sample/ack
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Sample/$exit
      -- CP-element group 334: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_sample_complete
      -- 
    ack_834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 334_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_offset_ack_0, ack => access_T_CP_0_elements(334)); -- 
    -- CP-element group 335:  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	331 
    -- CP-element group 335:  members (8) 
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_base_plus_offset/$entry
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_base_plus_offset/sum_rename_ack
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_base_plus_offset/sum_rename_req
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_base_plus_offset/$exit
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Update/ack
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_final_index_sum_regn_Update/$exit
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_offset_calculated
      -- CP-element group 335: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_137_root_address_calculated
      -- 
    ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_137_index_offset_ack_1, ack => access_T_CP_0_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	331 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	333 
    -- CP-element group 336: 	331 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_request/ack
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_request/$exit
      -- CP-element group 336: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_sample_completed_
      -- 
    ack_849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_138_final_reg_ack_0, ack => access_T_CP_0_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	332 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	338 
    -- CP-element group 337:  members (19) 
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_plus_offset/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_plus_offset/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_complete/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_addr_resize/base_resize_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_addr_resize/base_resize_req
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_addr_resize/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_addr_resize/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_address_resized
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_root_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_word_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_address_calculated
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_138_complete/ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_word_addrgen/root_register_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_word_addrgen/root_register_req
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_word_addrgen/$exit
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_word_addrgen/$entry
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_plus_offset/sum_rename_ack
      -- CP-element group 337: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_base_plus_offset/sum_rename_req
      -- 
    ack_854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_138_final_reg_ack_1, ack => access_T_CP_0_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	337 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (5) 
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_sample_start_
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/word_0/rr
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/word_0/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/$entry
      -- CP-element group 338: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/$entry
      -- 
    rr_887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(338), ack => ptr_deref_142_load_0_req_0); -- 
    access_T_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(337) & access_T_CP_0_elements(340);
      gj_access_T_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	347 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (5) 
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/word_0/cr
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_update_start_
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/word_0/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/$entry
      -- CP-element group 339: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/$entry
      -- 
    cr_898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(339), ack => ptr_deref_142_load_0_req_1); -- 
    access_T_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(347);
      gj_access_T_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: 	332 
    -- CP-element group 340:  members (5) 
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_sample_completed_
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/word_0/ra
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/word_0/$exit
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/word_access_start/$exit
      -- CP-element group 340: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Sample/$exit
      -- 
    ra_888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_142_load_0_ack_0, ack => access_T_CP_0_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	346 
    -- CP-element group 341:  members (9) 
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/ptr_deref_142_Merge/merge_ack
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/ptr_deref_142_Merge/merge_req
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/ptr_deref_142_Merge/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/ptr_deref_142_Merge/$entry
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_update_completed_
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/word_0/ca
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/word_0/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/word_access_complete/$exit
      -- CP-element group 341: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_142_Update/$exit
      -- 
    ca_899_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_142_load_0_ack_1, ack => access_T_CP_0_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	60 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Sample/req
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Sample/$entry
      -- CP-element group 342: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_sample_start_
      -- 
    req_912_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_912_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(342), ack => W_send_flag1_186_delayed_13_0_186_inst_req_0); -- 
    access_T_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(60) & access_T_CP_0_elements(344);
      gj_access_T_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	347 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Update/req
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_update_start_
      -- 
    req_917_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_917_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(343), ack => W_send_flag1_186_delayed_13_0_186_inst_req_1); -- 
    access_T_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(347);
      gj_access_T_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	56 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Sample/ack
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Sample/$exit
      -- CP-element group 344: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_sample_completed_
      -- 
    ack_913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag1_186_delayed_13_0_186_inst_ack_0, ack => access_T_CP_0_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	346 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Update/ack
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_188_update_completed_
      -- 
    ack_918_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag1_186_delayed_13_0_186_inst_ack_1, ack => access_T_CP_0_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	341 
    -- CP-element group 346: 	345 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	347 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_sample_start_
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Sample/req
      -- CP-element group 346: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Sample/$entry
      -- 
    req_926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(346), ack => WPIPE_input_pipe1_190_inst_req_0); -- 
    access_T_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(341) & access_T_CP_0_elements(345) & access_T_CP_0_elements(348);
      gj_access_T_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	346 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	348 
    -- CP-element group 347: marked-successors 
    -- CP-element group 347: 	339 
    -- CP-element group 347: 	343 
    -- CP-element group 347:  members (6) 
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_update_start_
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Update/req
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Sample/ack
      -- CP-element group 347: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Sample/$exit
      -- 
    ack_927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_190_inst_ack_0, ack => access_T_CP_0_elements(347)); -- 
    req_931_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_931_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(347), ack => WPIPE_input_pipe1_190_inst_req_1); -- 
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	347 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	404 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	346 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Update/ack
      -- CP-element group 348: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe1_190_Update/$exit
      -- 
    ack_932_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe1_190_inst_ack_1, ack => access_T_CP_0_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	353 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	354 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	354 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_request/req
      -- CP-element group 349: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_request/$entry
      -- 
    req_972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(349), ack => addr_of_204_final_reg_req_0); -- 
    access_T_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(353) & access_T_CP_0_elements(354);
      gj_access_T_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	9 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	358 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	355 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_complete/req
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_complete/$entry
      -- CP-element group 350: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_update_start_
      -- 
    req_977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(350), ack => addr_of_204_final_reg_req_1); -- 
    access_T_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(358);
      gj_access_T_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	9 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	354 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_update_start
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Update/req
      -- CP-element group 351: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Update/$entry
      -- 
    req_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(351), ack => array_obj_ref_203_index_offset_req_1); -- 
    access_T_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(354);
      gj_access_T_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	98 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	404 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	94 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Sample/ack
      -- CP-element group 352: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_sample_complete
      -- 
    ack_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_index_offset_ack_0, ack => access_T_CP_0_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	349 
    -- CP-element group 353:  members (8) 
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_base_plus_offset/$exit
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Update/ack
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_base_plus_offset/$entry
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_final_index_sum_regn_Update/$exit
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_offset_calculated
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_root_address_calculated
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_ack
      -- CP-element group 353: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_203_base_plus_offset/sum_rename_req
      -- 
    ack_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_203_index_offset_ack_1, ack => access_T_CP_0_elements(353)); -- 
    -- CP-element group 354:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: successors 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	349 
    -- CP-element group 354: 	351 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_request/ack
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_request/$exit
      -- CP-element group 354: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_sample_completed_
      -- 
    ack_973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 354_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_204_final_reg_ack_0, ack => access_T_CP_0_elements(354)); -- 
    -- CP-element group 355:  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	350 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	356 
    -- CP-element group 355:  members (19) 
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_complete/ack
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_complete/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_addr_resize/base_resize_ack
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_word_addrgen/root_register_ack
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_word_addrgen/root_register_req
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_word_addrgen/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_word_addrgen/$entry
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_plus_offset/sum_rename_ack
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_plus_offset/sum_rename_req
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_204_update_completed_
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_plus_offset/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_plus_offset/$entry
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_addr_resize/base_resize_req
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_addr_resize/$exit
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_addr_resize/$entry
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_address_resized
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_root_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_word_address_calculated
      -- CP-element group 355: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_base_address_calculated
      -- 
    ack_978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_204_final_reg_ack_1, ack => access_T_CP_0_elements(355)); -- 
    -- CP-element group 356:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	355 
    -- CP-element group 356: marked-predecessors 
    -- CP-element group 356: 	358 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	358 
    -- CP-element group 356:  members (5) 
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/$entry
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/word_0/rr
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/word_0/$entry
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/$entry
      -- CP-element group 356: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_sample_start_
      -- 
    rr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(356), ack => ptr_deref_208_load_0_req_0); -- 
    access_T_cp_element_group_356: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_356"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(355) & access_T_CP_0_elements(358);
      gj_access_T_cp_element_group_356 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(356), clk => clk, reset => reset); --
    end block;
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	365 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (5) 
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/$entry
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_update_start_
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/word_0/cr
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/word_0/$entry
      -- CP-element group 357: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/$entry
      -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(357), ack => ptr_deref_208_load_0_req_1); -- 
    access_T_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	356 
    -- CP-element group 358: successors 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	350 
    -- CP-element group 358: 	356 
    -- CP-element group 358:  members (5) 
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/$exit
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/word_0/ra
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/word_0/$exit
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Sample/word_access_start/$exit
      -- CP-element group 358: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_sample_completed_
      -- 
    ra_1012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 358_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_208_load_0_ack_0, ack => access_T_CP_0_elements(358)); -- 
    -- CP-element group 359:  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	364 
    -- CP-element group 359:  members (9) 
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/$exit
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/ptr_deref_208_Merge/merge_ack
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/ptr_deref_208_Merge/merge_req
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/ptr_deref_208_Merge/$exit
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_update_completed_
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/ptr_deref_208_Merge/$entry
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/word_0/ca
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/word_0/$exit
      -- CP-element group 359: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_208_Update/word_access_complete/$exit
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_208_load_0_ack_1, ack => access_T_CP_0_elements(359)); -- 
    -- CP-element group 360:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	140 
    -- CP-element group 360: marked-predecessors 
    -- CP-element group 360: 	362 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	362 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Sample/req
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_sample_start_
      -- CP-element group 360: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Sample/$entry
      -- 
    req_1036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(360), ack => W_send_flag2_249_delayed_13_0_252_inst_req_0); -- 
    access_T_cp_element_group_360: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_360"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(140) & access_T_CP_0_elements(362);
      gj_access_T_cp_element_group_360 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(360), clk => clk, reset => reset); --
    end block;
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	365 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_update_start_
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Update/req
      -- CP-element group 361: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Update/$entry
      -- 
    req_1041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(361), ack => W_send_flag2_249_delayed_13_0_252_inst_req_1); -- 
    access_T_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(365);
      gj_access_T_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: successors 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	360 
    -- CP-element group 362: 	136 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Sample/ack
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_sample_completed_
      -- CP-element group 362: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Sample/$exit
      -- 
    ack_1037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 362_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag2_249_delayed_13_0_252_inst_ack_0, ack => access_T_CP_0_elements(362)); -- 
    -- CP-element group 363:  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	364 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Update/ack
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_Update/$exit
      -- CP-element group 363: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_254_update_completed_
      -- 
    ack_1042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag2_249_delayed_13_0_252_inst_ack_1, ack => access_T_CP_0_elements(363)); -- 
    -- CP-element group 364:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	363 
    -- CP-element group 364: 	359 
    -- CP-element group 364: marked-predecessors 
    -- CP-element group 364: 	366 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	365 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_sample_start_
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Sample/req
      -- CP-element group 364: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Sample/$entry
      -- 
    req_1050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(364), ack => WPIPE_input_pipe2_256_inst_req_0); -- 
    access_T_cp_element_group_364: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_364"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(363) & access_T_CP_0_elements(359) & access_T_CP_0_elements(366);
      gj_access_T_cp_element_group_364 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(364), clk => clk, reset => reset); --
    end block;
    -- CP-element group 365:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	364 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	366 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	361 
    -- CP-element group 365: 	357 
    -- CP-element group 365:  members (6) 
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_update_start_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Update/req
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_sample_completed_
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Update/$entry
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Sample/ack
      -- CP-element group 365: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Sample/$exit
      -- 
    ack_1051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_256_inst_ack_0, ack => access_T_CP_0_elements(365)); -- 
    req_1055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(365), ack => WPIPE_input_pipe2_256_inst_req_1); -- 
    -- CP-element group 366:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	365 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	404 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	364 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Update/ack
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_update_completed_
      -- CP-element group 366: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe2_256_Update/$exit
      -- 
    ack_1056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 366_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe2_256_inst_ack_1, ack => access_T_CP_0_elements(366)); -- 
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	371 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	372 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	372 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_sample_start_
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_request/$entry
      -- CP-element group 367: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_request/req
      -- 
    req_1096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(367), ack => addr_of_270_final_reg_req_0); -- 
    access_T_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(371) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	9 
    -- CP-element group 368: marked-predecessors 
    -- CP-element group 368: 	376 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	373 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_update_start_
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_complete/$entry
      -- CP-element group 368: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_complete/req
      -- 
    req_1101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(368), ack => addr_of_270_final_reg_req_1); -- 
    access_T_cp_element_group_368: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_368"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(376);
      gj_access_T_cp_element_group_368 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(368), clk => clk, reset => reset); --
    end block;
    -- CP-element group 369:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	9 
    -- CP-element group 369: marked-predecessors 
    -- CP-element group 369: 	372 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Update/$entry
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Update/req
      -- CP-element group 369: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_update_start
      -- 
    req_1086_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1086_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(369), ack => array_obj_ref_269_index_offset_req_1); -- 
    access_T_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(372);
      gj_access_T_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	178 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	404 
    -- CP-element group 370: marked-successors 
    -- CP-element group 370: 	174 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/ack
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Sample/$exit
      -- CP-element group 370: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_sample_complete
      -- 
    ack_1082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 370_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_index_offset_ack_0, ack => access_T_CP_0_elements(370)); -- 
    -- CP-element group 371:  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	367 
    -- CP-element group 371:  members (8) 
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_root_address_calculated
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_offset_calculated
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Update/$exit
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_final_index_sum_regn_Update/ack
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_base_plus_offset/$entry
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_base_plus_offset/$exit
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_base_plus_offset/sum_rename_req
      -- CP-element group 371: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_269_base_plus_offset/sum_rename_ack
      -- 
    ack_1087_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_index_offset_ack_1, ack => access_T_CP_0_elements(371)); -- 
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	367 
    -- CP-element group 372: successors 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	367 
    -- CP-element group 372: 	369 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_request/$exit
      -- CP-element group 372: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_request/ack
      -- 
    ack_1097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_270_final_reg_ack_0, ack => access_T_CP_0_elements(372)); -- 
    -- CP-element group 373:  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	368 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (19) 
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_complete/$exit
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_270_complete/ack
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_address_calculated
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_word_address_calculated
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_root_address_calculated
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_address_resized
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_addr_resize/$entry
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_addr_resize/$exit
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_addr_resize/base_resize_req
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_addr_resize/base_resize_ack
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_plus_offset/$entry
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_plus_offset/$exit
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_plus_offset/sum_rename_req
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_base_plus_offset/sum_rename_ack
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_word_addrgen/$entry
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_word_addrgen/$exit
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_word_addrgen/root_register_req
      -- CP-element group 373: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_word_addrgen/root_register_ack
      -- 
    ack_1102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_270_final_reg_ack_1, ack => access_T_CP_0_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	373 
    -- CP-element group 374: marked-predecessors 
    -- CP-element group 374: 	376 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (5) 
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/$entry
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/word_0/$entry
      -- CP-element group 374: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/word_0/rr
      -- 
    rr_1135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(374), ack => ptr_deref_274_load_0_req_0); -- 
    access_T_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(373) & access_T_CP_0_elements(376);
      gj_access_T_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	383 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (5) 
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_update_start_
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/$entry
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/word_0/$entry
      -- CP-element group 375: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/word_0/cr
      -- 
    cr_1146_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1146_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(375), ack => ptr_deref_274_load_0_req_1); -- 
    access_T_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(383);
      gj_access_T_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: marked-successors 
    -- CP-element group 376: 	368 
    -- CP-element group 376: 	374 
    -- CP-element group 376:  members (5) 
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/$exit
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/word_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Sample/word_access_start/word_0/ra
      -- 
    ra_1136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_274_load_0_ack_0, ack => access_T_CP_0_elements(376)); -- 
    -- CP-element group 377:  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	382 
    -- CP-element group 377:  members (9) 
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/$exit
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/word_0/$exit
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/word_access_complete/word_0/ca
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/ptr_deref_274_Merge/$entry
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/ptr_deref_274_Merge/$exit
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/ptr_deref_274_Merge/merge_req
      -- CP-element group 377: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_274_Update/ptr_deref_274_Merge/merge_ack
      -- 
    ca_1147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_274_load_0_ack_1, ack => access_T_CP_0_elements(377)); -- 
    -- CP-element group 378:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	220 
    -- CP-element group 378: marked-predecessors 
    -- CP-element group 378: 	380 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Sample/req
      -- 
    req_1160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(378), ack => W_send_flag3_312_delayed_13_0_318_inst_req_0); -- 
    access_T_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(220) & access_T_CP_0_elements(380);
      gj_access_T_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	383 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_update_start_
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Update/req
      -- 
    req_1165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(379), ack => W_send_flag3_312_delayed_13_0_318_inst_req_1); -- 
    access_T_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(383);
      gj_access_T_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: marked-successors 
    -- CP-element group 380: 	216 
    -- CP-element group 380: 	378 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Sample/ack
      -- 
    ack_1161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag3_312_delayed_13_0_318_inst_ack_0, ack => access_T_CP_0_elements(380)); -- 
    -- CP-element group 381:  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	382 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_320_Update/ack
      -- 
    ack_1166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag3_312_delayed_13_0_318_inst_ack_1, ack => access_T_CP_0_elements(381)); -- 
    -- CP-element group 382:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	377 
    -- CP-element group 382: 	381 
    -- CP-element group 382: marked-predecessors 
    -- CP-element group 382: 	384 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	383 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_sample_start_
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Sample/$entry
      -- CP-element group 382: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Sample/req
      -- 
    req_1174_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1174_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(382), ack => WPIPE_input_pipe3_322_inst_req_0); -- 
    access_T_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(377) & access_T_CP_0_elements(381) & access_T_CP_0_elements(384);
      gj_access_T_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	382 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	384 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	375 
    -- CP-element group 383: 	379 
    -- CP-element group 383:  members (6) 
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_update_start_
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Sample/ack
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Update/$entry
      -- CP-element group 383: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Update/req
      -- 
    ack_1175_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_322_inst_ack_0, ack => access_T_CP_0_elements(383)); -- 
    req_1179_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1179_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(383), ack => WPIPE_input_pipe3_322_inst_req_1); -- 
    -- CP-element group 384:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	383 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	404 
    -- CP-element group 384: marked-successors 
    -- CP-element group 384: 	382 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe3_322_Update/ack
      -- 
    ack_1180_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe3_322_inst_ack_1, ack => access_T_CP_0_elements(384)); -- 
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	389 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	390 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	390 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_request/$entry
      -- CP-element group 385: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_request/req
      -- 
    req_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(385), ack => addr_of_336_final_reg_req_0); -- 
    access_T_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(389) & access_T_CP_0_elements(390);
      gj_access_T_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	9 
    -- CP-element group 386: marked-predecessors 
    -- CP-element group 386: 	394 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	391 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_update_start_
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_complete/$entry
      -- CP-element group 386: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_complete/req
      -- 
    req_1225_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1225_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(386), ack => addr_of_336_final_reg_req_1); -- 
    access_T_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(394);
      gj_access_T_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	9 
    -- CP-element group 387: marked-predecessors 
    -- CP-element group 387: 	390 
    -- CP-element group 387: successors 
    -- CP-element group 387: 	389 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_update_start
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Update/$entry
      -- CP-element group 387: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Update/req
      -- 
    req_1210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(387), ack => array_obj_ref_335_index_offset_req_1); -- 
    access_T_cp_element_group_387: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_387"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(9) & access_T_CP_0_elements(390);
      gj_access_T_cp_element_group_387 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(387), clk => clk, reset => reset); --
    end block;
    -- CP-element group 388:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	258 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	404 
    -- CP-element group 388: marked-successors 
    -- CP-element group 388: 	254 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_sample_complete
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Sample/$exit
      -- CP-element group 388: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Sample/ack
      -- 
    ack_1206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_335_index_offset_ack_0, ack => access_T_CP_0_elements(388)); -- 
    -- CP-element group 389:  transition  input  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	387 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	385 
    -- CP-element group 389:  members (8) 
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_root_address_calculated
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_offset_calculated
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Update/$exit
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_final_index_sum_regn_Update/ack
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_base_plus_offset/$entry
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_base_plus_offset/$exit
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_base_plus_offset/sum_rename_req
      -- CP-element group 389: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/array_obj_ref_335_base_plus_offset/sum_rename_ack
      -- 
    ack_1211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 389_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_335_index_offset_ack_1, ack => access_T_CP_0_elements(389)); -- 
    -- CP-element group 390:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	385 
    -- CP-element group 390: successors 
    -- CP-element group 390: marked-successors 
    -- CP-element group 390: 	385 
    -- CP-element group 390: 	387 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_request/$exit
      -- CP-element group 390: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_request/ack
      -- 
    ack_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_336_final_reg_ack_0, ack => access_T_CP_0_elements(390)); -- 
    -- CP-element group 391:  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	386 
    -- CP-element group 391: successors 
    -- CP-element group 391: 	392 
    -- CP-element group 391:  members (19) 
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_complete/$exit
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/addr_of_336_complete/ack
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_word_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_root_address_calculated
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_address_resized
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_addr_resize/$entry
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_addr_resize/$exit
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_addr_resize/base_resize_req
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_addr_resize/base_resize_ack
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_plus_offset/$entry
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_plus_offset/$exit
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_plus_offset/sum_rename_req
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_base_plus_offset/sum_rename_ack
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_word_addrgen/$entry
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_word_addrgen/$exit
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_word_addrgen/root_register_req
      -- CP-element group 391: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_word_addrgen/root_register_ack
      -- 
    ack_1226_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_336_final_reg_ack_1, ack => access_T_CP_0_elements(391)); -- 
    -- CP-element group 392:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	391 
    -- CP-element group 392: marked-predecessors 
    -- CP-element group 392: 	394 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	394 
    -- CP-element group 392:  members (5) 
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_sample_start_
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/word_0/$entry
      -- CP-element group 392: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/word_0/rr
      -- 
    rr_1259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(392), ack => ptr_deref_340_load_0_req_0); -- 
    access_T_cp_element_group_392: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_392"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(391) & access_T_CP_0_elements(394);
      gj_access_T_cp_element_group_392 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(392), clk => clk, reset => reset); --
    end block;
    -- CP-element group 393:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: marked-predecessors 
    -- CP-element group 393: 	401 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (5) 
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_update_start_
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/word_0/$entry
      -- CP-element group 393: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/word_0/cr
      -- 
    cr_1270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(393), ack => ptr_deref_340_load_0_req_1); -- 
    access_T_cp_element_group_393: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_393"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(401);
      gj_access_T_cp_element_group_393 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 394:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	392 
    -- CP-element group 394: successors 
    -- CP-element group 394: marked-successors 
    -- CP-element group 394: 	386 
    -- CP-element group 394: 	392 
    -- CP-element group 394:  members (5) 
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_sample_completed_
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/$exit
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/$exit
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/word_0/$exit
      -- CP-element group 394: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Sample/word_access_start/word_0/ra
      -- 
    ra_1260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 394_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_340_load_0_ack_0, ack => access_T_CP_0_elements(394)); -- 
    -- CP-element group 395:  transition  input  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: successors 
    -- CP-element group 395: 	400 
    -- CP-element group 395:  members (9) 
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_update_completed_
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/word_0/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/word_access_complete/word_0/ca
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/ptr_deref_340_Merge/$entry
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/ptr_deref_340_Merge/$exit
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/ptr_deref_340_Merge/merge_req
      -- CP-element group 395: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/ptr_deref_340_Update/ptr_deref_340_Merge/merge_ack
      -- 
    ca_1271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_340_load_0_ack_1, ack => access_T_CP_0_elements(395)); -- 
    -- CP-element group 396:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	300 
    -- CP-element group 396: marked-predecessors 
    -- CP-element group 396: 	398 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	398 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_sample_start_
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Sample/$entry
      -- CP-element group 396: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Sample/req
      -- 
    req_1284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(396), ack => W_send_flag4_375_delayed_13_0_384_inst_req_0); -- 
    access_T_cp_element_group_396: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_396"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= access_T_CP_0_elements(300) & access_T_CP_0_elements(398);
      gj_access_T_cp_element_group_396 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(396), clk => clk, reset => reset); --
    end block;
    -- CP-element group 397:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: marked-predecessors 
    -- CP-element group 397: 	401 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_update_start_
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Update/$entry
      -- CP-element group 397: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Update/req
      -- 
    req_1289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(397), ack => W_send_flag4_375_delayed_13_0_384_inst_req_1); -- 
    access_T_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= access_T_CP_0_elements(401);
      gj_access_T_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: successors 
    -- CP-element group 398: marked-successors 
    -- CP-element group 398: 	396 
    -- CP-element group 398: 	296 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_sample_completed_
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Sample/$exit
      -- CP-element group 398: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Sample/ack
      -- 
    ack_1285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 398_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag4_375_delayed_13_0_384_inst_ack_0, ack => access_T_CP_0_elements(398)); -- 
    -- CP-element group 399:  transition  input  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399: 	400 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_update_completed_
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Update/$exit
      -- CP-element group 399: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/assign_stmt_386_Update/ack
      -- 
    ack_1290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_flag4_375_delayed_13_0_384_inst_ack_1, ack => access_T_CP_0_elements(399)); -- 
    -- CP-element group 400:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	395 
    -- CP-element group 400: 	399 
    -- CP-element group 400: marked-predecessors 
    -- CP-element group 400: 	402 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	401 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_sample_start_
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Sample/$entry
      -- CP-element group 400: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Sample/req
      -- 
    req_1298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(400), ack => WPIPE_input_pipe4_388_inst_req_0); -- 
    access_T_cp_element_group_400: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_400"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= access_T_CP_0_elements(395) & access_T_CP_0_elements(399) & access_T_CP_0_elements(402);
      gj_access_T_cp_element_group_400 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(400), clk => clk, reset => reset); --
    end block;
    -- CP-element group 401:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	400 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	402 
    -- CP-element group 401: marked-successors 
    -- CP-element group 401: 	393 
    -- CP-element group 401: 	397 
    -- CP-element group 401:  members (6) 
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_sample_completed_
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_update_start_
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Sample/$exit
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Sample/ack
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Update/$entry
      -- CP-element group 401: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Update/req
      -- 
    ack_1299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 401_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_388_inst_ack_0, ack => access_T_CP_0_elements(401)); -- 
    req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => access_T_CP_0_elements(401), ack => WPIPE_input_pipe4_388_inst_req_1); -- 
    -- CP-element group 402:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	401 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402: marked-successors 
    -- CP-element group 402: 	400 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_update_completed_
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Update/$exit
      -- CP-element group 402: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/WPIPE_input_pipe4_388_Update/ack
      -- 
    ack_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 402_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_pipe4_388_inst_ack_1, ack => access_T_CP_0_elements(402)); -- 
    -- CP-element group 403:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	9 
    -- CP-element group 403: successors 
    -- CP-element group 403: 	10 
    -- CP-element group 403:  members (1) 
      -- CP-element group 403: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group access_T_CP_0_elements(403) is a control-delay.
    cp_element_403_delay: control_delay_element  generic map(name => " 403_delay", delay_value => 1)  port map(req => access_T_CP_0_elements(9), ack => access_T_CP_0_elements(403), clk => clk, reset =>reset);
    -- CP-element group 404:  join  transition  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	334 
    -- CP-element group 404: 	366 
    -- CP-element group 404: 	370 
    -- CP-element group 404: 	384 
    -- CP-element group 404: 	388 
    -- CP-element group 404: 	402 
    -- CP-element group 404: 	12 
    -- CP-element group 404: 	348 
    -- CP-element group 404: 	352 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	6 
    -- CP-element group 404:  members (1) 
      -- CP-element group 404: 	 branch_block_stmt_29/do_while_stmt_42/do_while_stmt_42_loop_body/$exit
      -- 
    access_T_cp_element_group_404: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 29) := "access_T_cp_element_group_404"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= access_T_CP_0_elements(334) & access_T_CP_0_elements(366) & access_T_CP_0_elements(370) & access_T_CP_0_elements(384) & access_T_CP_0_elements(388) & access_T_CP_0_elements(402) & access_T_CP_0_elements(12) & access_T_CP_0_elements(348) & access_T_CP_0_elements(352);
      gj_access_T_cp_element_group_404 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => access_T_CP_0_elements(404), clk => clk, reset => reset); --
    end block;
    -- CP-element group 405:  transition  input  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	5 
    -- CP-element group 405: successors 
    -- CP-element group 405:  members (2) 
      -- CP-element group 405: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/$exit
      -- CP-element group 405: 	 branch_block_stmt_29/do_while_stmt_42/loop_exit/ack
      -- 
    ack_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 405_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_42_branch_ack_0, ack => access_T_CP_0_elements(405)); -- 
    -- CP-element group 406:  transition  input  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	5 
    -- CP-element group 406: successors 
    -- CP-element group 406:  members (2) 
      -- CP-element group 406: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/$exit
      -- CP-element group 406: 	 branch_block_stmt_29/do_while_stmt_42/loop_taken/ack
      -- 
    ack_1313_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 406_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_42_branch_ack_1, ack => access_T_CP_0_elements(406)); -- 
    -- CP-element group 407:  transition  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	3 
    -- CP-element group 407: successors 
    -- CP-element group 407: 	1 
    -- CP-element group 407:  members (1) 
      -- CP-element group 407: 	 branch_block_stmt_29/do_while_stmt_42/$exit
      -- 
    access_T_CP_0_elements(407) <= access_T_CP_0_elements(3);
    access_T_do_while_stmt_42_terminator_1314: loop_terminator -- 
      generic map (name => " access_T_do_while_stmt_42_terminator_1314", max_iterations_in_flight =>15) 
      port map(loop_body_exit => access_T_CP_0_elements(6),loop_continue => access_T_CP_0_elements(406),loop_terminate => access_T_CP_0_elements(405),loop_back => access_T_CP_0_elements(4),loop_exit => access_T_CP_0_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_44_phi_seq_78_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(23);
      access_T_CP_0_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(26);
      access_T_CP_0_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(28);
      access_T_CP_0_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(21);
      access_T_CP_0_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(32);
      access_T_CP_0_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(33);
      access_T_CP_0_elements(22) <= phi_mux_reqs(1);
      phi_stmt_44_phi_seq_78 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_44_phi_seq_78") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(17), 
          phi_sample_ack => access_T_CP_0_elements(18), 
          phi_update_req => access_T_CP_0_elements(19), 
          phi_update_ack => access_T_CP_0_elements(20), 
          phi_mux_ack => access_T_CP_0_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_49_phi_seq_132_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(42);
      access_T_CP_0_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(49);
      access_T_CP_0_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(50);
      access_T_CP_0_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(40);
      access_T_CP_0_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(53);
      access_T_CP_0_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(54);
      access_T_CP_0_elements(41) <= phi_mux_reqs(1);
      phi_stmt_49_phi_seq_132 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_49_phi_seq_132") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(36), 
          phi_sample_ack => access_T_CP_0_elements(37), 
          phi_update_req => access_T_CP_0_elements(38), 
          phi_update_ack => access_T_CP_0_elements(39), 
          phi_mux_ack => access_T_CP_0_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_54_phi_seq_176_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(63);
      access_T_CP_0_elements(66)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(66);
      access_T_CP_0_elements(67)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(68);
      access_T_CP_0_elements(64) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(61);
      access_T_CP_0_elements(70)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(72);
      access_T_CP_0_elements(71)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(73);
      access_T_CP_0_elements(62) <= phi_mux_reqs(1);
      phi_stmt_54_phi_seq_176 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_54_phi_seq_176") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(57), 
          phi_sample_ack => access_T_CP_0_elements(58), 
          phi_update_req => access_T_CP_0_elements(59), 
          phi_update_ack => access_T_CP_0_elements(60), 
          phi_mux_ack => access_T_CP_0_elements(65), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_59_phi_seq_220_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(80);
      access_T_CP_0_elements(85)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(87);
      access_T_CP_0_elements(86)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(88);
      access_T_CP_0_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(82);
      access_T_CP_0_elements(89)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(89);
      access_T_CP_0_elements(90)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(91);
      access_T_CP_0_elements(83) <= phi_mux_reqs(1);
      phi_stmt_59_phi_seq_220 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_59_phi_seq_220") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(76), 
          phi_sample_ack => access_T_CP_0_elements(77), 
          phi_update_req => access_T_CP_0_elements(78), 
          phi_update_ack => access_T_CP_0_elements(79), 
          phi_mux_ack => access_T_CP_0_elements(84), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_64_phi_seq_274_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(99);
      access_T_CP_0_elements(104)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(106);
      access_T_CP_0_elements(105)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(107);
      access_T_CP_0_elements(100) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(101);
      access_T_CP_0_elements(108)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(112);
      access_T_CP_0_elements(109)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(113);
      access_T_CP_0_elements(102) <= phi_mux_reqs(1);
      phi_stmt_64_phi_seq_274 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_64_phi_seq_274") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(95), 
          phi_sample_ack => access_T_CP_0_elements(96), 
          phi_update_req => access_T_CP_0_elements(97), 
          phi_update_ack => access_T_CP_0_elements(98), 
          phi_mux_ack => access_T_CP_0_elements(103), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_69_phi_seq_328_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(120);
      access_T_CP_0_elements(125)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(127);
      access_T_CP_0_elements(126)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(128);
      access_T_CP_0_elements(121) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(122);
      access_T_CP_0_elements(129)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(133);
      access_T_CP_0_elements(130)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(134);
      access_T_CP_0_elements(123) <= phi_mux_reqs(1);
      phi_stmt_69_phi_seq_328 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_69_phi_seq_328") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(116), 
          phi_sample_ack => access_T_CP_0_elements(117), 
          phi_update_req => access_T_CP_0_elements(118), 
          phi_update_ack => access_T_CP_0_elements(119), 
          phi_mux_ack => access_T_CP_0_elements(124), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_74_phi_seq_372_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(143);
      access_T_CP_0_elements(146)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(146);
      access_T_CP_0_elements(147)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(148);
      access_T_CP_0_elements(144) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(141);
      access_T_CP_0_elements(150)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(152);
      access_T_CP_0_elements(151)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(153);
      access_T_CP_0_elements(142) <= phi_mux_reqs(1);
      phi_stmt_74_phi_seq_372 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_74_phi_seq_372") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(137), 
          phi_sample_ack => access_T_CP_0_elements(138), 
          phi_update_req => access_T_CP_0_elements(139), 
          phi_update_ack => access_T_CP_0_elements(140), 
          phi_mux_ack => access_T_CP_0_elements(145), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_79_phi_seq_416_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(162);
      access_T_CP_0_elements(165)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(165);
      access_T_CP_0_elements(166)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(167);
      access_T_CP_0_elements(163) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(160);
      access_T_CP_0_elements(169)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(171);
      access_T_CP_0_elements(170)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(172);
      access_T_CP_0_elements(161) <= phi_mux_reqs(1);
      phi_stmt_79_phi_seq_416 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_79_phi_seq_416") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(156), 
          phi_sample_ack => access_T_CP_0_elements(157), 
          phi_update_req => access_T_CP_0_elements(158), 
          phi_update_ack => access_T_CP_0_elements(159), 
          phi_mux_ack => access_T_CP_0_elements(164), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_84_phi_seq_470_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(179);
      access_T_CP_0_elements(184)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(186);
      access_T_CP_0_elements(185)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(187);
      access_T_CP_0_elements(180) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(181);
      access_T_CP_0_elements(188)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(192);
      access_T_CP_0_elements(189)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(193);
      access_T_CP_0_elements(182) <= phi_mux_reqs(1);
      phi_stmt_84_phi_seq_470 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_84_phi_seq_470") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(175), 
          phi_sample_ack => access_T_CP_0_elements(176), 
          phi_update_req => access_T_CP_0_elements(177), 
          phi_update_ack => access_T_CP_0_elements(178), 
          phi_mux_ack => access_T_CP_0_elements(183), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_89_phi_seq_524_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(200);
      access_T_CP_0_elements(205)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(207);
      access_T_CP_0_elements(206)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(208);
      access_T_CP_0_elements(201) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(202);
      access_T_CP_0_elements(209)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(213);
      access_T_CP_0_elements(210)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(214);
      access_T_CP_0_elements(203) <= phi_mux_reqs(1);
      phi_stmt_89_phi_seq_524 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_89_phi_seq_524") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(196), 
          phi_sample_ack => access_T_CP_0_elements(197), 
          phi_update_req => access_T_CP_0_elements(198), 
          phi_update_ack => access_T_CP_0_elements(199), 
          phi_mux_ack => access_T_CP_0_elements(204), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_94_phi_seq_568_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(223);
      access_T_CP_0_elements(226)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(226);
      access_T_CP_0_elements(227)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(228);
      access_T_CP_0_elements(224) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(221);
      access_T_CP_0_elements(230)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(232);
      access_T_CP_0_elements(231)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(233);
      access_T_CP_0_elements(222) <= phi_mux_reqs(1);
      phi_stmt_94_phi_seq_568 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_94_phi_seq_568") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(217), 
          phi_sample_ack => access_T_CP_0_elements(218), 
          phi_update_req => access_T_CP_0_elements(219), 
          phi_update_ack => access_T_CP_0_elements(220), 
          phi_mux_ack => access_T_CP_0_elements(225), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_99_phi_seq_612_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(240);
      access_T_CP_0_elements(245)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(247);
      access_T_CP_0_elements(246)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(248);
      access_T_CP_0_elements(241) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(242);
      access_T_CP_0_elements(249)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(249);
      access_T_CP_0_elements(250)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(251);
      access_T_CP_0_elements(243) <= phi_mux_reqs(1);
      phi_stmt_99_phi_seq_612 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_99_phi_seq_612") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(236), 
          phi_sample_ack => access_T_CP_0_elements(237), 
          phi_update_req => access_T_CP_0_elements(238), 
          phi_update_ack => access_T_CP_0_elements(239), 
          phi_mux_ack => access_T_CP_0_elements(244), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_104_phi_seq_666_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(261);
      access_T_CP_0_elements(264)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(268);
      access_T_CP_0_elements(265)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(269);
      access_T_CP_0_elements(262) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(259);
      access_T_CP_0_elements(270)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(272);
      access_T_CP_0_elements(271)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(273);
      access_T_CP_0_elements(260) <= phi_mux_reqs(1);
      phi_stmt_104_phi_seq_666 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_104_phi_seq_666") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(255), 
          phi_sample_ack => access_T_CP_0_elements(256), 
          phi_update_req => access_T_CP_0_elements(257), 
          phi_update_ack => access_T_CP_0_elements(258), 
          phi_mux_ack => access_T_CP_0_elements(263), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_111_phi_seq_720_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(280);
      access_T_CP_0_elements(285)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(287);
      access_T_CP_0_elements(286)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(288);
      access_T_CP_0_elements(281) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(282);
      access_T_CP_0_elements(289)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(293);
      access_T_CP_0_elements(290)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(294);
      access_T_CP_0_elements(283) <= phi_mux_reqs(1);
      phi_stmt_111_phi_seq_720 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_111_phi_seq_720") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(276), 
          phi_sample_ack => access_T_CP_0_elements(277), 
          phi_update_req => access_T_CP_0_elements(278), 
          phi_update_ack => access_T_CP_0_elements(279), 
          phi_mux_ack => access_T_CP_0_elements(284), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_116_phi_seq_764_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(303);
      access_T_CP_0_elements(306)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(306);
      access_T_CP_0_elements(307)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(308);
      access_T_CP_0_elements(304) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(301);
      access_T_CP_0_elements(310)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(312);
      access_T_CP_0_elements(311)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(313);
      access_T_CP_0_elements(302) <= phi_mux_reqs(1);
      phi_stmt_116_phi_seq_764 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_116_phi_seq_764") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(297), 
          phi_sample_ack => access_T_CP_0_elements(298), 
          phi_update_req => access_T_CP_0_elements(299), 
          phi_update_ack => access_T_CP_0_elements(300), 
          phi_mux_ack => access_T_CP_0_elements(305), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_121_phi_seq_808_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= access_T_CP_0_elements(318);
      access_T_CP_0_elements(323)<= src_sample_reqs(0);
      src_sample_acks(0)  <= access_T_CP_0_elements(325);
      access_T_CP_0_elements(324)<= src_update_reqs(0);
      src_update_acks(0)  <= access_T_CP_0_elements(326);
      access_T_CP_0_elements(319) <= phi_mux_reqs(0);
      triggers(1)  <= access_T_CP_0_elements(320);
      access_T_CP_0_elements(327)<= src_sample_reqs(1);
      src_sample_acks(1)  <= access_T_CP_0_elements(327);
      access_T_CP_0_elements(328)<= src_update_reqs(1);
      src_update_acks(1)  <= access_T_CP_0_elements(329);
      access_T_CP_0_elements(321) <= phi_mux_reqs(1);
      phi_stmt_121_phi_seq_808 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_121_phi_seq_808") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => access_T_CP_0_elements(11), 
          phi_sample_ack => access_T_CP_0_elements(316), 
          phi_update_req => access_T_CP_0_elements(13), 
          phi_update_ack => access_T_CP_0_elements(317), 
          phi_mux_ack => access_T_CP_0_elements(322), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= access_T_CP_0_elements(7);
        preds(1)  <= access_T_CP_0_elements(8);
        entry_tmerge_30 : transition_merge -- 
          generic map(name => " entry_tmerge_30")
          port map (preds => preds, symbol_out => access_T_CP_0_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_162_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_228_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_294_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_360_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_108_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_171_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_237_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_303_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_369_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_34_wire : std_logic_vector(15 downto 0);
    signal MUX_173_wire : std_logic_vector(31 downto 0);
    signal MUX_239_wire : std_logic_vector(31 downto 0);
    signal MUX_305_wire : std_logic_vector(31 downto 0);
    signal MUX_371_wire : std_logic_vector(31 downto 0);
    signal OR_u1_u1_394_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_397_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_398_wire : std_logic_vector(0 downto 0);
    signal address1_44 : std_logic_vector(31 downto 0);
    signal address2_64 : std_logic_vector(31 downto 0);
    signal address3_84 : std_logic_vector(31 downto 0);
    signal address4_104 : std_logic_vector(31 downto 0);
    signal array_obj_ref_137_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_137_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_137_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_137_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_137_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_137_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_203_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_269_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_335_root_address : std_logic_vector(13 downto 0);
    signal continue_flag1_185 : std_logic_vector(0 downto 0);
    signal continue_flag2_251 : std_logic_vector(0 downto 0);
    signal continue_flag3_317 : std_logic_vector(0 downto 0);
    signal continue_flag4_383 : std_logic_vector(0 downto 0);
    signal fetch_addr1_139 : std_logic_vector(31 downto 0);
    signal fetch_addr2_205 : std_logic_vector(31 downto 0);
    signal fetch_addr3_271 : std_logic_vector(31 downto 0);
    signal fetch_addr4_337 : std_logic_vector(31 downto 0);
    signal fv1_143 : std_logic_vector(63 downto 0);
    signal fv2_209 : std_logic_vector(63 downto 0);
    signal fv3_275 : std_logic_vector(63 downto 0);
    signal fv4_341 : std_logic_vector(63 downto 0);
    signal konst_129_wire_constant : std_logic_vector(31 downto 0);
    signal konst_149_wire_constant : std_logic_vector(31 downto 0);
    signal konst_161_wire_constant : std_logic_vector(15 downto 0);
    signal konst_172_wire_constant : std_logic_vector(31 downto 0);
    signal konst_195_wire_constant : std_logic_vector(31 downto 0);
    signal konst_215_wire_constant : std_logic_vector(31 downto 0);
    signal konst_227_wire_constant : std_logic_vector(15 downto 0);
    signal konst_238_wire_constant : std_logic_vector(31 downto 0);
    signal konst_261_wire_constant : std_logic_vector(31 downto 0);
    signal konst_281_wire_constant : std_logic_vector(31 downto 0);
    signal konst_293_wire_constant : std_logic_vector(15 downto 0);
    signal konst_304_wire_constant : std_logic_vector(31 downto 0);
    signal konst_327_wire_constant : std_logic_vector(31 downto 0);
    signal konst_347_wire_constant : std_logic_vector(31 downto 0);
    signal konst_359_wire_constant : std_logic_vector(15 downto 0);
    signal konst_370_wire_constant : std_logic_vector(31 downto 0);
    signal konst_39_wire_constant : std_logic_vector(31 downto 0);
    signal m2_factor_41 : std_logic_vector(31 downto 0);
    signal m_factor_36 : std_logic_vector(31 downto 0);
    signal mycounter1_49 : std_logic_vector(31 downto 0);
    signal mycounter2_69 : std_logic_vector(31 downto 0);
    signal mycounter3_89 : std_logic_vector(31 downto 0);
    signal mycounter4_111 : std_logic_vector(31 downto 0);
    signal n_address1_175 : std_logic_vector(31 downto 0);
    signal n_address1_175_48_buffered : std_logic_vector(31 downto 0);
    signal n_address2_241 : std_logic_vector(31 downto 0);
    signal n_address2_241_66_buffered : std_logic_vector(31 downto 0);
    signal n_address3_307 : std_logic_vector(31 downto 0);
    signal n_address3_307_86_buffered : std_logic_vector(31 downto 0);
    signal n_address4_373 : std_logic_vector(31 downto 0);
    signal n_address4_373_110_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter1_157 : std_logic_vector(31 downto 0);
    signal n_mycounter1_157_53_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter2_223 : std_logic_vector(31 downto 0);
    signal n_mycounter2_223_71_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter3_289 : std_logic_vector(31 downto 0);
    signal n_mycounter3_289_91_buffered : std_logic_vector(31 downto 0);
    signal n_mycounter4_355 : std_logic_vector(31 downto 0);
    signal n_mycounter4_355_113_buffered : std_logic_vector(31 downto 0);
    signal n_row1_165 : std_logic_vector(15 downto 0);
    signal n_row1_165_58_buffered : std_logic_vector(15 downto 0);
    signal n_row2_231 : std_logic_vector(15 downto 0);
    signal n_row2_231_78_buffered : std_logic_vector(15 downto 0);
    signal n_row3_297 : std_logic_vector(15 downto 0);
    signal n_row3_297_98_buffered : std_logic_vector(15 downto 0);
    signal n_row4_363 : std_logic_vector(15 downto 0);
    signal n_row4_363_120_buffered : std_logic_vector(15 downto 0);
    signal n_start1_146 : std_logic_vector(0 downto 0);
    signal n_start1_146_61_buffered : std_logic_vector(0 downto 0);
    signal n_start2_212 : std_logic_vector(0 downto 0);
    signal n_start2_212_83_buffered : std_logic_vector(0 downto 0);
    signal n_start3_278 : std_logic_vector(0 downto 0);
    signal n_start3_278_101_buffered : std_logic_vector(0 downto 0);
    signal n_start4_344 : std_logic_vector(0 downto 0);
    signal n_start4_344_123_buffered : std_logic_vector(0 downto 0);
    signal next_row1_131 : std_logic_vector(0 downto 0);
    signal next_row2_197 : std_logic_vector(0 downto 0);
    signal next_row3_263 : std_logic_vector(0 downto 0);
    signal next_row4_329 : std_logic_vector(0 downto 0);
    signal ptr_deref_142_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_142_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_142_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_142_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_142_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_208_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_208_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_208_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_208_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_208_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_274_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_274_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_274_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_274_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_274_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_340_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_340_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_340_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_340_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_340_word_offset_0 : std_logic_vector(13 downto 0);
    signal row1_54 : std_logic_vector(15 downto 0);
    signal row2_74 : std_logic_vector(15 downto 0);
    signal row3_94 : std_logic_vector(15 downto 0);
    signal row4_116 : std_logic_vector(15 downto 0);
    signal send_flag1_180 : std_logic_vector(0 downto 0);
    signal send_flag1_186_delayed_13_0_188 : std_logic_vector(0 downto 0);
    signal send_flag2_246 : std_logic_vector(0 downto 0);
    signal send_flag2_249_delayed_13_0_254 : std_logic_vector(0 downto 0);
    signal send_flag3_312 : std_logic_vector(0 downto 0);
    signal send_flag3_312_delayed_13_0_320 : std_logic_vector(0 downto 0);
    signal send_flag4_375_delayed_13_0_386 : std_logic_vector(0 downto 0);
    signal send_flag4_378 : std_logic_vector(0 downto 0);
    signal start1_59 : std_logic_vector(0 downto 0);
    signal start2_79 : std_logic_vector(0 downto 0);
    signal start3_99 : std_logic_vector(0 downto 0);
    signal start4_121 : std_logic_vector(0 downto 0);
    signal tmp_cnt1_151 : std_logic_vector(31 downto 0);
    signal tmp_cnt2_217 : std_logic_vector(31 downto 0);
    signal tmp_cnt3_283 : std_logic_vector(31 downto 0);
    signal tmp_cnt4_349 : std_logic_vector(31 downto 0);
    signal type_cast_103_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_109_wire : std_logic_vector(31 downto 0);
    signal type_cast_115_wire : std_logic_vector(31 downto 0);
    signal type_cast_119_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_125_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_136_resized : std_logic_vector(13 downto 0);
    signal type_cast_136_scaled : std_logic_vector(13 downto 0);
    signal type_cast_136_wire : std_logic_vector(63 downto 0);
    signal type_cast_202_resized : std_logic_vector(13 downto 0);
    signal type_cast_202_scaled : std_logic_vector(13 downto 0);
    signal type_cast_202_wire : std_logic_vector(63 downto 0);
    signal type_cast_268_resized : std_logic_vector(13 downto 0);
    signal type_cast_268_scaled : std_logic_vector(13 downto 0);
    signal type_cast_268_wire : std_logic_vector(63 downto 0);
    signal type_cast_334_resized : std_logic_vector(13 downto 0);
    signal type_cast_334_scaled : std_logic_vector(13 downto 0);
    signal type_cast_334_wire : std_logic_vector(63 downto 0);
    signal type_cast_47_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_52_wire : std_logic_vector(31 downto 0);
    signal type_cast_57_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_63_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_68_wire : std_logic_vector(31 downto 0);
    signal type_cast_73_wire : std_logic_vector(31 downto 0);
    signal type_cast_77_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_82_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_88_wire : std_logic_vector(31 downto 0);
    signal type_cast_93_wire : std_logic_vector(31 downto 0);
    signal type_cast_97_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_137_constant_part_of_offset <= "00000000000000";
    array_obj_ref_137_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_137_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_137_resized_base_address <= "00000000000000";
    array_obj_ref_203_constant_part_of_offset <= "00000000000000";
    array_obj_ref_203_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_203_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_203_resized_base_address <= "00000000000000";
    array_obj_ref_269_constant_part_of_offset <= "00000000000000";
    array_obj_ref_269_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_269_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_269_resized_base_address <= "00000000000000";
    array_obj_ref_335_constant_part_of_offset <= "00000000000000";
    array_obj_ref_335_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_335_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_335_resized_base_address <= "00000000000000";
    konst_129_wire_constant <= "00000000000000000000000000000001";
    konst_149_wire_constant <= "00000000000000000000000000000001";
    konst_161_wire_constant <= "0000000000000010";
    konst_172_wire_constant <= "00000000000000000000000000000001";
    konst_195_wire_constant <= "00000000000000000000000000000001";
    konst_215_wire_constant <= "00000000000000000000000000000001";
    konst_227_wire_constant <= "0000000000000010";
    konst_238_wire_constant <= "00000000000000000000000000000001";
    konst_261_wire_constant <= "00000000000000000000000000000001";
    konst_281_wire_constant <= "00000000000000000000000000000001";
    konst_293_wire_constant <= "0000000000000010";
    konst_304_wire_constant <= "00000000000000000000000000000001";
    konst_327_wire_constant <= "00000000000000000000000000000001";
    konst_347_wire_constant <= "00000000000000000000000000000001";
    konst_359_wire_constant <= "0000000000000010";
    konst_370_wire_constant <= "00000000000000000000000000000001";
    konst_39_wire_constant <= "00000000000000000000000000000001";
    ptr_deref_142_word_offset_0 <= "00000000000000";
    ptr_deref_208_word_offset_0 <= "00000000000000";
    ptr_deref_274_word_offset_0 <= "00000000000000";
    ptr_deref_340_word_offset_0 <= "00000000000000";
    type_cast_103_wire_constant <= "1";
    type_cast_119_wire_constant <= "0000000000000001";
    type_cast_125_wire_constant <= "1";
    type_cast_47_wire_constant <= "00000000000000000000000000000000";
    type_cast_57_wire_constant <= "0000000000000000";
    type_cast_63_wire_constant <= "1";
    type_cast_77_wire_constant <= "0000000000000000";
    type_cast_82_wire_constant <= "1";
    type_cast_97_wire_constant <= "0000000000000000";
    phi_stmt_104: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_109_wire & n_address4_373_110_buffered;
      req <= phi_stmt_104_req_0 & phi_stmt_104_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_104",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_104_ack_0,
          idata => idata,
          odata => address4_104,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_104
    phi_stmt_111: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_mycounter4_355_113_buffered & type_cast_115_wire;
      req <= phi_stmt_111_req_0 & phi_stmt_111_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_111",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_111_ack_0,
          idata => idata,
          odata => mycounter4_111,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_111
    phi_stmt_116: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_119_wire_constant & n_row4_363_120_buffered;
      req <= phi_stmt_116_req_0 & phi_stmt_116_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_116",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_116_ack_0,
          idata => idata,
          odata => row4_116,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_116
    phi_stmt_121: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_start4_344_123_buffered & type_cast_125_wire_constant;
      req <= phi_stmt_121_req_0 & phi_stmt_121_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_121",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_121_ack_0,
          idata => idata,
          odata => start4_121,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_121
    phi_stmt_44: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_47_wire_constant & n_address1_175_48_buffered;
      req <= phi_stmt_44_req_0 & phi_stmt_44_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_44",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_44_ack_0,
          idata => idata,
          odata => address1_44,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_44
    phi_stmt_49: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_52_wire & n_mycounter1_157_53_buffered;
      req <= phi_stmt_49_req_0 & phi_stmt_49_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_49",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_49_ack_0,
          idata => idata,
          odata => mycounter1_49,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_49
    phi_stmt_54: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_57_wire_constant & n_row1_165_58_buffered;
      req <= phi_stmt_54_req_0 & phi_stmt_54_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_54",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_54_ack_0,
          idata => idata,
          odata => row1_54,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_54
    phi_stmt_59: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_start1_146_61_buffered & type_cast_63_wire_constant;
      req <= phi_stmt_59_req_0 & phi_stmt_59_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_59",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_59_ack_0,
          idata => idata,
          odata => start1_59,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_59
    phi_stmt_64: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address2_241_66_buffered & type_cast_68_wire;
      req <= phi_stmt_64_req_0 & phi_stmt_64_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_64",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_64_ack_0,
          idata => idata,
          odata => address2_64,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_64
    phi_stmt_69: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_mycounter2_223_71_buffered & type_cast_73_wire;
      req <= phi_stmt_69_req_0 & phi_stmt_69_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_69",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_69_ack_0,
          idata => idata,
          odata => mycounter2_69,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_69
    phi_stmt_74: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_77_wire_constant & n_row2_231_78_buffered;
      req <= phi_stmt_74_req_0 & phi_stmt_74_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_74",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_74_ack_0,
          idata => idata,
          odata => row2_74,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_74
    phi_stmt_79: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_82_wire_constant & n_start2_212_83_buffered;
      req <= phi_stmt_79_req_0 & phi_stmt_79_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_79",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_79_ack_0,
          idata => idata,
          odata => start2_79,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_79
    phi_stmt_84: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_address3_307_86_buffered & type_cast_88_wire;
      req <= phi_stmt_84_req_0 & phi_stmt_84_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_84",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_84_ack_0,
          idata => idata,
          odata => address3_84,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_84
    phi_stmt_89: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_mycounter3_289_91_buffered & type_cast_93_wire;
      req <= phi_stmt_89_req_0 & phi_stmt_89_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_89",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_89_ack_0,
          idata => idata,
          odata => mycounter3_89,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_89
    phi_stmt_94: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_97_wire_constant & n_row3_297_98_buffered;
      req <= phi_stmt_94_req_0 & phi_stmt_94_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_94",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_94_ack_0,
          idata => idata,
          odata => row3_94,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_94
    phi_stmt_99: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_start3_278_101_buffered & type_cast_103_wire_constant;
      req <= phi_stmt_99_req_0 & phi_stmt_99_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_99",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_99_ack_0,
          idata => idata,
          odata => start3_99,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_99
    -- flow-through select operator MUX_156_inst
    n_mycounter1_157 <= m_factor_36 when (next_row1_131(0) /=  '0') else tmp_cnt1_151;
    -- flow-through select operator MUX_164_inst
    n_row1_165 <= ADD_u16_u16_162_wire when (next_row1_131(0) /=  '0') else row1_54;
    -- flow-through select operator MUX_173_inst
    MUX_173_wire <= ADD_u32_u32_171_wire when (next_row1_131(0) /=  '0') else konst_172_wire_constant;
    -- flow-through select operator MUX_222_inst
    n_mycounter2_223 <= m_factor_36 when (next_row2_197(0) /=  '0') else tmp_cnt2_217;
    -- flow-through select operator MUX_230_inst
    n_row2_231 <= ADD_u16_u16_228_wire when (next_row2_197(0) /=  '0') else row2_74;
    -- flow-through select operator MUX_239_inst
    MUX_239_wire <= ADD_u32_u32_237_wire when (next_row2_197(0) /=  '0') else konst_238_wire_constant;
    -- flow-through select operator MUX_288_inst
    n_mycounter3_289 <= m_factor_36 when (next_row3_263(0) /=  '0') else tmp_cnt3_283;
    -- flow-through select operator MUX_296_inst
    n_row3_297 <= ADD_u16_u16_294_wire when (next_row3_263(0) /=  '0') else row3_94;
    -- flow-through select operator MUX_305_inst
    MUX_305_wire <= ADD_u32_u32_303_wire when (next_row3_263(0) /=  '0') else konst_304_wire_constant;
    -- flow-through select operator MUX_354_inst
    n_mycounter4_355 <= m_factor_36 when (next_row4_329(0) /=  '0') else tmp_cnt4_349;
    -- flow-through select operator MUX_362_inst
    n_row4_363 <= ADD_u16_u16_360_wire when (next_row4_329(0) /=  '0') else row4_116;
    -- flow-through select operator MUX_371_inst
    MUX_371_wire <= ADD_u32_u32_369_wire when (next_row4_329(0) /=  '0') else konst_370_wire_constant;
    -- interlock W_n_start1_144_inst
    process(next_row1_131) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row1_131(0 downto 0);
      n_start1_146 <= tmp_var; -- 
    end process;
    -- interlock W_n_start2_210_inst
    process(next_row2_197) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row2_197(0 downto 0);
      n_start2_212 <= tmp_var; -- 
    end process;
    -- interlock W_n_start3_276_inst
    process(next_row3_263) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row3_263(0 downto 0);
      n_start3_278 <= tmp_var; -- 
    end process;
    -- interlock W_n_start4_342_inst
    process(next_row4_329) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := next_row4_329(0 downto 0);
      n_start4_344 <= tmp_var; -- 
    end process;
    W_send_flag1_186_delayed_13_0_186_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_flag1_186_delayed_13_0_186_inst_req_0;
      W_send_flag1_186_delayed_13_0_186_inst_ack_0<= wack(0);
      rreq(0) <= W_send_flag1_186_delayed_13_0_186_inst_req_1;
      W_send_flag1_186_delayed_13_0_186_inst_ack_1<= rack(0);
      W_send_flag1_186_delayed_13_0_186_inst : InterlockBuffer generic map ( -- 
        name => "W_send_flag1_186_delayed_13_0_186_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_flag1_180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_flag1_186_delayed_13_0_188,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_flag2_249_delayed_13_0_252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_flag2_249_delayed_13_0_252_inst_req_0;
      W_send_flag2_249_delayed_13_0_252_inst_ack_0<= wack(0);
      rreq(0) <= W_send_flag2_249_delayed_13_0_252_inst_req_1;
      W_send_flag2_249_delayed_13_0_252_inst_ack_1<= rack(0);
      W_send_flag2_249_delayed_13_0_252_inst : InterlockBuffer generic map ( -- 
        name => "W_send_flag2_249_delayed_13_0_252_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_flag2_246,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_flag2_249_delayed_13_0_254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_flag3_312_delayed_13_0_318_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_flag3_312_delayed_13_0_318_inst_req_0;
      W_send_flag3_312_delayed_13_0_318_inst_ack_0<= wack(0);
      rreq(0) <= W_send_flag3_312_delayed_13_0_318_inst_req_1;
      W_send_flag3_312_delayed_13_0_318_inst_ack_1<= rack(0);
      W_send_flag3_312_delayed_13_0_318_inst : InterlockBuffer generic map ( -- 
        name => "W_send_flag3_312_delayed_13_0_318_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_flag3_312,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_flag3_312_delayed_13_0_320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_flag4_375_delayed_13_0_384_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_flag4_375_delayed_13_0_384_inst_req_0;
      W_send_flag4_375_delayed_13_0_384_inst_ack_0<= wack(0);
      rreq(0) <= W_send_flag4_375_delayed_13_0_384_inst_req_1;
      W_send_flag4_375_delayed_13_0_384_inst_ack_1<= rack(0);
      W_send_flag4_375_delayed_13_0_384_inst : InterlockBuffer generic map ( -- 
        name => "W_send_flag4_375_delayed_13_0_384_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_flag4_378,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_flag4_375_delayed_13_0_386,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_138_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_138_final_reg_req_0;
      addr_of_138_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_138_final_reg_req_1;
      addr_of_138_final_reg_ack_1<= rack(0);
      addr_of_138_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_138_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_137_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_204_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_204_final_reg_req_0;
      addr_of_204_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_204_final_reg_req_1;
      addr_of_204_final_reg_ack_1<= rack(0);
      addr_of_204_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_204_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_203_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_205,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_270_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_270_final_reg_req_0;
      addr_of_270_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_270_final_reg_req_1;
      addr_of_270_final_reg_ack_1<= rack(0);
      addr_of_270_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_270_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_269_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr3_271,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_336_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_336_final_reg_req_0;
      addr_of_336_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_336_final_reg_req_1;
      addr_of_336_final_reg_ack_1<= rack(0);
      addr_of_336_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_336_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_335_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr4_337,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_175_48_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_175_48_buf_req_0;
      n_address1_175_48_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_175_48_buf_req_1;
      n_address1_175_48_buf_ack_1<= rack(0);
      n_address1_175_48_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_175_48_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_175,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_175_48_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_241_66_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_241_66_buf_req_0;
      n_address2_241_66_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_241_66_buf_req_1;
      n_address2_241_66_buf_ack_1<= rack(0);
      n_address2_241_66_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_241_66_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_241_66_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address3_307_86_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address3_307_86_buf_req_0;
      n_address3_307_86_buf_ack_0<= wack(0);
      rreq(0) <= n_address3_307_86_buf_req_1;
      n_address3_307_86_buf_ack_1<= rack(0);
      n_address3_307_86_buf : InterlockBuffer generic map ( -- 
        name => "n_address3_307_86_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address3_307,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address3_307_86_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address4_373_110_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address4_373_110_buf_req_0;
      n_address4_373_110_buf_ack_0<= wack(0);
      rreq(0) <= n_address4_373_110_buf_req_1;
      n_address4_373_110_buf_ack_1<= rack(0);
      n_address4_373_110_buf : InterlockBuffer generic map ( -- 
        name => "n_address4_373_110_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address4_373,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address4_373_110_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter1_157_53_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter1_157_53_buf_req_0;
      n_mycounter1_157_53_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter1_157_53_buf_req_1;
      n_mycounter1_157_53_buf_ack_1<= rack(0);
      n_mycounter1_157_53_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter1_157_53_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter1_157,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter1_157_53_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter2_223_71_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter2_223_71_buf_req_0;
      n_mycounter2_223_71_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter2_223_71_buf_req_1;
      n_mycounter2_223_71_buf_ack_1<= rack(0);
      n_mycounter2_223_71_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter2_223_71_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter2_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter2_223_71_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter3_289_91_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter3_289_91_buf_req_0;
      n_mycounter3_289_91_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter3_289_91_buf_req_1;
      n_mycounter3_289_91_buf_ack_1<= rack(0);
      n_mycounter3_289_91_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter3_289_91_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter3_289,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter3_289_91_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_mycounter4_355_113_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_mycounter4_355_113_buf_req_0;
      n_mycounter4_355_113_buf_ack_0<= wack(0);
      rreq(0) <= n_mycounter4_355_113_buf_req_1;
      n_mycounter4_355_113_buf_ack_1<= rack(0);
      n_mycounter4_355_113_buf : InterlockBuffer generic map ( -- 
        name => "n_mycounter4_355_113_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_mycounter4_355,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_mycounter4_355_113_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row1_165_58_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row1_165_58_buf_req_0;
      n_row1_165_58_buf_ack_0<= wack(0);
      rreq(0) <= n_row1_165_58_buf_req_1;
      n_row1_165_58_buf_ack_1<= rack(0);
      n_row1_165_58_buf : InterlockBuffer generic map ( -- 
        name => "n_row1_165_58_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row1_165,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row1_165_58_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row2_231_78_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row2_231_78_buf_req_0;
      n_row2_231_78_buf_ack_0<= wack(0);
      rreq(0) <= n_row2_231_78_buf_req_1;
      n_row2_231_78_buf_ack_1<= rack(0);
      n_row2_231_78_buf : InterlockBuffer generic map ( -- 
        name => "n_row2_231_78_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row2_231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row2_231_78_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row3_297_98_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row3_297_98_buf_req_0;
      n_row3_297_98_buf_ack_0<= wack(0);
      rreq(0) <= n_row3_297_98_buf_req_1;
      n_row3_297_98_buf_ack_1<= rack(0);
      n_row3_297_98_buf : InterlockBuffer generic map ( -- 
        name => "n_row3_297_98_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row3_297,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row3_297_98_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row4_363_120_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row4_363_120_buf_req_0;
      n_row4_363_120_buf_ack_0<= wack(0);
      rreq(0) <= n_row4_363_120_buf_req_1;
      n_row4_363_120_buf_ack_1<= rack(0);
      n_row4_363_120_buf : InterlockBuffer generic map ( -- 
        name => "n_row4_363_120_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row4_363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row4_363_120_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start1_146_61_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start1_146_61_buf_req_0;
      n_start1_146_61_buf_ack_0<= wack(0);
      rreq(0) <= n_start1_146_61_buf_req_1;
      n_start1_146_61_buf_ack_1<= rack(0);
      n_start1_146_61_buf : InterlockBuffer generic map ( -- 
        name => "n_start1_146_61_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start1_146,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start1_146_61_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start2_212_83_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start2_212_83_buf_req_0;
      n_start2_212_83_buf_ack_0<= wack(0);
      rreq(0) <= n_start2_212_83_buf_req_1;
      n_start2_212_83_buf_ack_1<= rack(0);
      n_start2_212_83_buf : InterlockBuffer generic map ( -- 
        name => "n_start2_212_83_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start2_212,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start2_212_83_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start3_278_101_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start3_278_101_buf_req_0;
      n_start3_278_101_buf_ack_0<= wack(0);
      rreq(0) <= n_start3_278_101_buf_req_1;
      n_start3_278_101_buf_ack_1<= rack(0);
      n_start3_278_101_buf : InterlockBuffer generic map ( -- 
        name => "n_start3_278_101_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start3_278,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start3_278_101_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_start4_344_123_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_start4_344_123_buf_req_0;
      n_start4_344_123_buf_ack_0<= wack(0);
      rreq(0) <= n_start4_344_123_buf_req_1;
      n_start4_344_123_buf_ack_1<= rack(0);
      n_start4_344_123_buf : InterlockBuffer generic map ( -- 
        name => "n_start4_344_123_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_start4_344,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_start4_344_123_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_109_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_109_inst_req_0;
      type_cast_109_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_109_inst_req_1;
      type_cast_109_inst_ack_1<= rack(0);
      type_cast_109_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_109_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ADD_u32_u32_108_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_109_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_115_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_115_inst_req_0;
      type_cast_115_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_115_inst_req_1;
      type_cast_115_inst_ack_1<= rack(0);
      type_cast_115_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_115_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_115_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_136_inst
    process(address1_44) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := address1_44(31 downto 0);
      type_cast_136_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_202_inst
    process(address2_64) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := address2_64(31 downto 0);
      type_cast_202_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_268_inst
    process(address3_84) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := address3_84(31 downto 0);
      type_cast_268_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_334_inst
    process(address4_104) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := address4_104(31 downto 0);
      type_cast_334_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_35_inst
    process(MUL_u16_u16_34_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_34_wire(15 downto 0);
      m_factor_36 <= tmp_var; -- 
    end process;
    type_cast_52_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_52_inst_req_0;
      type_cast_52_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_52_inst_req_1;
      type_cast_52_inst_ack_1<= rack(0);
      type_cast_52_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_52_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_52_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_68_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_68_inst_req_0;
      type_cast_68_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_68_inst_req_1;
      type_cast_68_inst_ack_1<= rack(0);
      type_cast_68_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_68_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_68_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_73_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_73_inst_req_0;
      type_cast_73_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_73_inst_req_1;
      type_cast_73_inst_ack_1<= rack(0);
      type_cast_73_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_73_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_73_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_88_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_88_inst_req_0;
      type_cast_88_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_88_inst_req_1;
      type_cast_88_inst_ack_1<= rack(0);
      type_cast_88_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_88_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m2_factor_41,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_88_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_93_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_93_inst_req_0;
      type_cast_93_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_93_inst_req_1;
      type_cast_93_inst_ack_1<= rack(0);
      type_cast_93_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_93_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => m_factor_36,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_93_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_137_index_1_rename
    process(type_cast_136_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_136_resized;
      ov(13 downto 0) := iv;
      type_cast_136_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_index_1_resize
    process(type_cast_136_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_136_wire;
      ov := iv(13 downto 0);
      type_cast_136_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_137_root_address_inst
    process(array_obj_ref_137_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_137_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_137_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_1_rename
    process(type_cast_202_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_202_resized;
      ov(13 downto 0) := iv;
      type_cast_202_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_index_1_resize
    process(type_cast_202_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_202_wire;
      ov := iv(13 downto 0);
      type_cast_202_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_203_root_address_inst
    process(array_obj_ref_203_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_203_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_203_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_index_1_rename
    process(type_cast_268_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_268_resized;
      ov(13 downto 0) := iv;
      type_cast_268_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_index_1_resize
    process(type_cast_268_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_268_wire;
      ov := iv(13 downto 0);
      type_cast_268_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_269_root_address_inst
    process(array_obj_ref_269_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_269_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_269_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_index_1_rename
    process(type_cast_334_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_334_resized;
      ov(13 downto 0) := iv;
      type_cast_334_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_index_1_resize
    process(type_cast_334_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_334_wire;
      ov := iv(13 downto 0);
      type_cast_334_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_335_root_address_inst
    process(array_obj_ref_335_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_335_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_335_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_addr_0
    process(ptr_deref_142_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_142_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_base_resize
    process(fetch_addr1_139) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_139;
      ov := iv(13 downto 0);
      ptr_deref_142_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_gather_scatter
    process(ptr_deref_142_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_data_0;
      ov(63 downto 0) := iv;
      fv1_143 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_142_root_address_inst
    process(ptr_deref_142_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_142_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_142_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_208_addr_0
    process(ptr_deref_208_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_208_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_208_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_208_base_resize
    process(fetch_addr2_205) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_205;
      ov := iv(13 downto 0);
      ptr_deref_208_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_208_gather_scatter
    process(ptr_deref_208_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_208_data_0;
      ov(63 downto 0) := iv;
      fv2_209 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_208_root_address_inst
    process(ptr_deref_208_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_208_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_208_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_274_addr_0
    process(ptr_deref_274_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_274_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_274_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_274_base_resize
    process(fetch_addr3_271) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr3_271;
      ov := iv(13 downto 0);
      ptr_deref_274_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_274_gather_scatter
    process(ptr_deref_274_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_274_data_0;
      ov(63 downto 0) := iv;
      fv3_275 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_274_root_address_inst
    process(ptr_deref_274_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_274_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_274_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_addr_0
    process(ptr_deref_340_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_340_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_base_resize
    process(fetch_addr4_337) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr4_337;
      ov := iv(13 downto 0);
      ptr_deref_340_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_gather_scatter
    process(ptr_deref_340_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_data_0;
      ov(63 downto 0) := iv;
      fv4_341 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_340_root_address_inst
    process(ptr_deref_340_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_340_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_340_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_42_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= OR_u1_u1_398_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_42_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_42_branch_req_0,
          ack0 => do_while_stmt_42_branch_ack_0,
          ack1 => do_while_stmt_42_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_162_inst
    process(row1_54) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row1_54, konst_161_wire_constant, tmp_var);
      ADD_u16_u16_162_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_228_inst
    process(row2_74) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row2_74, konst_227_wire_constant, tmp_var);
      ADD_u16_u16_228_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_294_inst
    process(row3_94) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row3_94, konst_293_wire_constant, tmp_var);
      ADD_u16_u16_294_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_360_inst
    process(row4_116) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row4_116, konst_359_wire_constant, tmp_var);
      ADD_u16_u16_360_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_108_inst
    process(m_factor_36, m2_factor_41) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, m2_factor_41, tmp_var);
      ADD_u32_u32_108_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_171_inst
    process(m_factor_36, mycounter1_49) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter1_49, tmp_var);
      ADD_u32_u32_171_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_174_inst
    process(address1_44, MUX_173_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_44, MUX_173_wire, tmp_var);
      n_address1_175 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_237_inst
    process(m_factor_36, mycounter2_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter2_69, tmp_var);
      ADD_u32_u32_237_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_240_inst
    process(address2_64, MUX_239_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_64, MUX_239_wire, tmp_var);
      n_address2_241 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_303_inst
    process(m_factor_36, mycounter3_89) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter3_89, tmp_var);
      ADD_u32_u32_303_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_306_inst
    process(address3_84, MUX_305_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address3_84, MUX_305_wire, tmp_var);
      n_address3_307 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_369_inst
    process(m_factor_36, mycounter4_111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(m_factor_36, mycounter4_111, tmp_var);
      ADD_u32_u32_369_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_372_inst
    process(address4_104, MUX_371_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address4_104, MUX_371_wire, tmp_var);
      n_address4_373 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_130_inst
    process(mycounter1_49) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter1_49, konst_129_wire_constant, tmp_var);
      next_row1_131 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_196_inst
    process(mycounter2_69) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter2_69, konst_195_wire_constant, tmp_var);
      next_row2_197 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_262_inst
    process(mycounter3_89) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter3_89, konst_261_wire_constant, tmp_var);
      next_row3_263 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_328_inst
    process(mycounter4_111) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(mycounter4_111, konst_327_wire_constant, tmp_var);
      next_row4_329 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_34_inst
    process(ct_buffer, chl_in_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(ct_buffer, chl_in_buffer, tmp_var);
      MUL_u16_u16_34_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_394_inst
    process(continue_flag1_185, continue_flag2_251) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(continue_flag1_185, continue_flag2_251, tmp_var);
      OR_u1_u1_394_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_397_inst
    process(continue_flag3_317, continue_flag4_383) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(continue_flag3_317, continue_flag4_383, tmp_var);
      OR_u1_u1_397_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_398_inst
    process(OR_u1_u1_394_wire, OR_u1_u1_397_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_394_wire, OR_u1_u1_397_wire, tmp_var);
      OR_u1_u1_398_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_40_inst
    process(m_factor_36) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(m_factor_36, konst_39_wire_constant, tmp_var);
      m2_factor_41 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_150_inst
    process(mycounter1_49) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter1_49, konst_149_wire_constant, tmp_var);
      tmp_cnt1_151 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_216_inst
    process(mycounter2_69) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter2_69, konst_215_wire_constant, tmp_var);
      tmp_cnt2_217 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_282_inst
    process(mycounter3_89) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter3_89, konst_281_wire_constant, tmp_var);
      tmp_cnt3_283 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_348_inst
    process(mycounter4_111) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(mycounter4_111, konst_347_wire_constant, tmp_var);
      tmp_cnt4_349 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_179_inst
    process(row1_54, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row1_54, row_in_buffer, tmp_var);
      send_flag1_180 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_184_inst
    process(n_row1_165, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row1_165, row_in_buffer, tmp_var);
      continue_flag1_185 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_245_inst
    process(row2_74, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row2_74, row_in_buffer, tmp_var);
      send_flag2_246 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_250_inst
    process(n_row2_231, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row2_231, row_in_buffer, tmp_var);
      continue_flag2_251 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_311_inst
    process(row3_94, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row3_94, row_in_buffer, tmp_var);
      send_flag3_312 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_316_inst
    process(n_row3_297, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row3_297, row_in_buffer, tmp_var);
      continue_flag3_317 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_377_inst
    process(row4_116, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(row4_116, row_in_buffer, tmp_var);
      send_flag4_378 <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_382_inst
    process(n_row4_363, row_in_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(n_row4_363, row_in_buffer, tmp_var);
      continue_flag4_383 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_137_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_136_scaled;
      array_obj_ref_137_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_137_index_offset_req_0;
      array_obj_ref_137_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_137_index_offset_req_1;
      array_obj_ref_137_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_203_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_202_scaled;
      array_obj_ref_203_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_203_index_offset_req_0;
      array_obj_ref_203_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_203_index_offset_req_1;
      array_obj_ref_203_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_269_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_268_scaled;
      array_obj_ref_269_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_269_index_offset_req_0;
      array_obj_ref_269_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_269_index_offset_req_1;
      array_obj_ref_269_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : array_obj_ref_335_index_offset 
    ApIntAdd_group_37: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_334_scaled;
      array_obj_ref_335_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_335_index_offset_req_0;
      array_obj_ref_335_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_335_index_offset_req_1;
      array_obj_ref_335_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_37_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared load operator group (0) : ptr_deref_208_load_0 ptr_deref_142_load_0 ptr_deref_274_load_0 ptr_deref_340_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 6, 1 => 6, 2 => 6, 3 => 6);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_208_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_142_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_274_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_340_load_0_req_0;
      ptr_deref_208_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_142_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_274_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_340_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_208_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_142_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_274_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_340_load_0_req_1;
      ptr_deref_208_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_142_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_274_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_340_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 2) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 2) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_208_word_address_0 & ptr_deref_142_word_address_0 & ptr_deref_274_word_address_0 & ptr_deref_340_word_address_0;
      ptr_deref_208_data_0 <= data_out(255 downto 192);
      ptr_deref_142_data_0 <= data_out(191 downto 128);
      ptr_deref_274_data_0 <= data_out(127 downto 64);
      ptr_deref_340_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(13 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(63 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_input_pipe1_190_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe1_190_inst_req_0;
      WPIPE_input_pipe1_190_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe1_190_inst_req_1;
      WPIPE_input_pipe1_190_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag1_186_delayed_13_0_188(0);
      data_in <= fv1_143;
      input_pipe1_write_0_gI: SplitGuardInterface generic map(name => "input_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "input_pipe1", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe1_pipe_write_req(0),
          oack => input_pipe1_pipe_write_ack(0),
          odata => input_pipe1_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_input_pipe2_256_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe2_256_inst_req_0;
      WPIPE_input_pipe2_256_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe2_256_inst_req_1;
      WPIPE_input_pipe2_256_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag2_249_delayed_13_0_254(0);
      data_in <= fv2_209;
      input_pipe2_write_1_gI: SplitGuardInterface generic map(name => "input_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "input_pipe2", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe2_pipe_write_req(0),
          oack => input_pipe2_pipe_write_ack(0),
          odata => input_pipe2_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_input_pipe3_322_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe3_322_inst_req_0;
      WPIPE_input_pipe3_322_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe3_322_inst_req_1;
      WPIPE_input_pipe3_322_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag3_312_delayed_13_0_320(0);
      data_in <= fv3_275;
      input_pipe3_write_2_gI: SplitGuardInterface generic map(name => "input_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "input_pipe3", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe3_pipe_write_req(0),
          oack => input_pipe3_pipe_write_ack(0),
          odata => input_pipe3_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_input_pipe4_388_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_pipe4_388_inst_req_0;
      WPIPE_input_pipe4_388_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_pipe4_388_inst_req_1;
      WPIPE_input_pipe4_388_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_flag4_375_delayed_13_0_386(0);
      data_in <= fv4_341;
      input_pipe4_write_3_gI: SplitGuardInterface generic map(name => "input_pipe4_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_pipe4_write_3: OutputPortRevised -- 
        generic map ( name => "input_pipe4", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_pipe4_pipe_write_req(0),
          oack => input_pipe4_pipe_write_ack(0),
          odata => input_pipe4_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end access_T_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolution3D is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    timer_call_reqs : out  std_logic_vector(0 downto 0);
    timer_call_acks : in   std_logic_vector(0 downto 0);
    timer_call_tag  :  out  std_logic_vector(1 downto 0);
    timer_return_reqs : out  std_logic_vector(0 downto 0);
    timer_return_acks : in   std_logic_vector(0 downto 0);
    timer_return_data : in   std_logic_vector(63 downto 0);
    timer_return_tag :  in   std_logic_vector(1 downto 0);
    access_T_call_reqs : out  std_logic_vector(0 downto 0);
    access_T_call_acks : in   std_logic_vector(0 downto 0);
    access_T_call_data : out  std_logic_vector(47 downto 0);
    access_T_call_tag  :  out  std_logic_vector(0 downto 0);
    access_T_return_reqs : out  std_logic_vector(0 downto 0);
    access_T_return_acks : in   std_logic_vector(0 downto 0);
    access_T_return_tag :  in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_call_data : out  std_logic_vector(47 downto 0);
    loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
    loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
    loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
    sendB_call_reqs : out  std_logic_vector(0 downto 0);
    sendB_call_acks : in   std_logic_vector(0 downto 0);
    sendB_call_data : out  std_logic_vector(31 downto 0);
    sendB_call_tag  :  out  std_logic_vector(0 downto 0);
    sendB_return_reqs : out  std_logic_vector(0 downto 0);
    sendB_return_acks : in   std_logic_vector(0 downto 0);
    sendB_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolution3D;
architecture convolution3D_arch of convolution3D is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolution3D_CP_2151_start: Boolean;
  signal convolution3D_CP_2151_symbol: Boolean;
  -- volatile/operator module components. 
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(31 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal type_cast_739_inst_ack_0 : boolean;
  signal type_cast_739_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_797_inst_ack_0 : boolean;
  signal type_cast_814_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_735_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_735_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_722_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_785_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_772_inst_ack_1 : boolean;
  signal type_cast_764_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_1 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_785_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_785_inst_ack_0 : boolean;
  signal type_cast_801_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_772_inst_req_1 : boolean;
  signal type_cast_726_inst_ack_1 : boolean;
  signal type_cast_726_inst_req_1 : boolean;
  signal type_cast_789_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_747_inst_ack_1 : boolean;
  signal type_cast_789_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_747_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_860_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1402_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_860_inst_ack_1 : boolean;
  signal type_cast_751_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_860_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_860_inst_ack_0 : boolean;
  signal type_cast_851_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_835_inst_ack_0 : boolean;
  signal type_cast_851_inst_req_0 : boolean;
  signal type_cast_851_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1402_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_0 : boolean;
  signal type_cast_1334_inst_ack_1 : boolean;
  signal type_cast_839_inst_ack_1 : boolean;
  signal type_cast_1529_inst_req_1 : boolean;
  signal type_cast_839_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_req_0 : boolean;
  signal type_cast_826_inst_ack_0 : boolean;
  signal type_cast_826_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_835_inst_req_0 : boolean;
  signal type_cast_801_inst_req_0 : boolean;
  signal type_cast_1539_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1348_inst_req_0 : boolean;
  signal type_cast_826_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_797_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_822_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_822_inst_req_1 : boolean;
  signal type_cast_1462_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_822_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_822_inst_req_0 : boolean;
  signal if_stmt_1446_branch_ack_0 : boolean;
  signal type_cast_726_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_797_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_772_inst_ack_0 : boolean;
  signal type_cast_726_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_797_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_772_inst_req_0 : boolean;
  signal type_cast_851_inst_req_1 : boolean;
  signal type_cast_814_inst_ack_1 : boolean;
  signal type_cast_839_inst_ack_0 : boolean;
  signal type_cast_826_inst_ack_1 : boolean;
  signal type_cast_1334_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1348_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1348_inst_ack_1 : boolean;
  signal type_cast_1303_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_722_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_722_inst_req_1 : boolean;
  signal type_cast_801_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_735_inst_ack_1 : boolean;
  signal type_cast_764_inst_ack_1 : boolean;
  signal type_cast_801_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_735_inst_req_1 : boolean;
  signal type_cast_764_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_785_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_722_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_ack_0 : boolean;
  signal type_cast_864_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1402_inst_req_0 : boolean;
  signal type_cast_864_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_835_inst_ack_1 : boolean;
  signal type_cast_1462_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_835_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1299_inst_ack_0 : boolean;
  signal type_cast_776_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_885_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_885_inst_ack_1 : boolean;
  signal type_cast_1511_inst_ack_1 : boolean;
  signal array_obj_ref_1295_index_offset_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_810_inst_req_0 : boolean;
  signal type_cast_864_inst_req_1 : boolean;
  signal type_cast_889_inst_req_1 : boolean;
  signal type_cast_1388_inst_ack_1 : boolean;
  signal type_cast_889_inst_ack_1 : boolean;
  signal if_stmt_1563_branch_req_0 : boolean;
  signal type_cast_1511_inst_req_1 : boolean;
  signal type_cast_839_inst_req_0 : boolean;
  signal type_cast_1511_inst_req_0 : boolean;
  signal type_cast_889_inst_req_0 : boolean;
  signal type_cast_889_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_747_inst_ack_0 : boolean;
  signal type_cast_776_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1402_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_847_inst_ack_1 : boolean;
  signal type_cast_1334_inst_ack_0 : boolean;
  signal if_stmt_1446_branch_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1535_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_897_inst_req_0 : boolean;
  signal type_cast_1388_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_897_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_747_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_872_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_ack_0 : boolean;
  signal type_cast_1005_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_872_inst_req_1 : boolean;
  signal type_cast_776_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_760_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_872_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_872_inst_ack_0 : boolean;
  signal type_cast_776_inst_req_0 : boolean;
  signal if_stmt_1446_branch_ack_1 : boolean;
  signal type_cast_739_inst_ack_1 : boolean;
  signal type_cast_864_inst_ack_1 : boolean;
  signal type_cast_739_inst_req_1 : boolean;
  signal type_cast_1334_inst_req_1 : boolean;
  signal type_cast_814_inst_ack_0 : boolean;
  signal type_cast_876_inst_ack_1 : boolean;
  signal type_cast_814_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1348_inst_ack_0 : boolean;
  signal type_cast_789_inst_ack_1 : boolean;
  signal type_cast_1511_inst_ack_0 : boolean;
  signal type_cast_876_inst_req_1 : boolean;
  signal type_cast_789_inst_req_1 : boolean;
  signal type_cast_876_inst_req_0 : boolean;
  signal type_cast_876_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_885_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_885_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1299_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_ack_0 : boolean;
  signal type_cast_1303_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1299_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1299_inst_ack_1 : boolean;
  signal type_cast_1406_inst_req_0 : boolean;
  signal type_cast_764_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_897_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_897_inst_ack_1 : boolean;
  signal type_cast_901_inst_req_0 : boolean;
  signal type_cast_901_inst_ack_0 : boolean;
  signal type_cast_901_inst_req_1 : boolean;
  signal type_cast_901_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_910_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_910_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_910_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_910_inst_ack_1 : boolean;
  signal type_cast_914_inst_req_0 : boolean;
  signal type_cast_914_inst_ack_0 : boolean;
  signal type_cast_914_inst_req_1 : boolean;
  signal type_cast_914_inst_ack_1 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal type_cast_923_inst_req_1 : boolean;
  signal type_cast_923_inst_ack_1 : boolean;
  signal type_cast_927_inst_req_0 : boolean;
  signal type_cast_927_inst_ack_0 : boolean;
  signal type_cast_927_inst_req_1 : boolean;
  signal type_cast_927_inst_ack_1 : boolean;
  signal type_cast_1352_inst_ack_1 : boolean;
  signal array_obj_ref_1295_index_offset_req_0 : boolean;
  signal type_cast_1352_inst_req_1 : boolean;
  signal if_stmt_945_branch_req_0 : boolean;
  signal type_cast_1515_inst_req_1 : boolean;
  signal if_stmt_945_branch_ack_1 : boolean;
  signal if_stmt_945_branch_ack_0 : boolean;
  signal type_cast_1424_inst_ack_1 : boolean;
  signal type_cast_982_inst_req_0 : boolean;
  signal type_cast_982_inst_ack_0 : boolean;
  signal type_cast_1352_inst_ack_0 : boolean;
  signal type_cast_982_inst_req_1 : boolean;
  signal type_cast_982_inst_ack_1 : boolean;
  signal type_cast_1529_inst_ack_1 : boolean;
  signal if_stmt_1563_branch_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1535_inst_req_1 : boolean;
  signal type_cast_1424_inst_req_1 : boolean;
  signal ptr_deref_1432_store_0_ack_1 : boolean;
  signal type_cast_1424_inst_ack_0 : boolean;
  signal type_cast_1352_inst_req_0 : boolean;
  signal ptr_deref_1432_store_0_req_1 : boolean;
  signal array_obj_ref_1011_index_offset_req_0 : boolean;
  signal array_obj_ref_1011_index_offset_ack_0 : boolean;
  signal array_obj_ref_1011_index_offset_req_1 : boolean;
  signal type_cast_1388_inst_ack_0 : boolean;
  signal array_obj_ref_1011_index_offset_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1535_inst_ack_0 : boolean;
  signal type_cast_1388_inst_req_0 : boolean;
  signal addr_of_1012_final_reg_req_0 : boolean;
  signal addr_of_1012_final_reg_ack_0 : boolean;
  signal addr_of_1012_final_reg_req_1 : boolean;
  signal addr_of_1012_final_reg_ack_1 : boolean;
  signal type_cast_1424_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1015_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1015_inst_ack_0 : boolean;
  signal addr_of_1296_final_reg_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1535_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1015_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1015_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_req_1 : boolean;
  signal type_cast_1515_inst_ack_0 : boolean;
  signal type_cast_1019_inst_req_0 : boolean;
  signal type_cast_1019_inst_ack_0 : boolean;
  signal type_cast_1019_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_1 : boolean;
  signal type_cast_1019_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1028_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1028_inst_ack_0 : boolean;
  signal addr_of_1296_final_reg_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1028_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1028_inst_ack_1 : boolean;
  signal type_cast_1515_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_ack_0 : boolean;
  signal type_cast_1032_inst_req_0 : boolean;
  signal type_cast_1032_inst_ack_0 : boolean;
  signal type_cast_1032_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_ack_0 : boolean;
  signal type_cast_1032_inst_ack_1 : boolean;
  signal type_cast_1539_inst_ack_1 : boolean;
  signal ptr_deref_1432_store_0_ack_0 : boolean;
  signal ptr_deref_1432_store_0_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1046_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1384_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1046_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1046_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1046_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1330_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1420_inst_ack_1 : boolean;
  signal type_cast_1050_inst_req_0 : boolean;
  signal type_cast_1050_inst_ack_0 : boolean;
  signal type_cast_1050_inst_req_1 : boolean;
  signal type_cast_1050_inst_ack_1 : boolean;
  signal type_cast_1539_inst_req_1 : boolean;
  signal if_stmt_1563_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1852_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1420_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1064_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1064_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1064_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1064_inst_ack_1 : boolean;
  signal type_cast_1068_inst_req_0 : boolean;
  signal type_cast_1068_inst_ack_0 : boolean;
  signal type_cast_1068_inst_req_1 : boolean;
  signal type_cast_1068_inst_ack_1 : boolean;
  signal addr_of_1296_final_reg_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1082_inst_req_0 : boolean;
  signal type_cast_1370_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1082_inst_ack_0 : boolean;
  signal addr_of_1296_final_reg_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1082_inst_req_1 : boolean;
  signal type_cast_1370_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1082_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1420_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1420_inst_req_0 : boolean;
  signal if_stmt_1486_branch_ack_0 : boolean;
  signal type_cast_1086_inst_req_0 : boolean;
  signal type_cast_1086_inst_ack_0 : boolean;
  signal type_cast_1086_inst_req_1 : boolean;
  signal type_cast_1086_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1100_inst_req_0 : boolean;
  signal type_cast_1370_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1100_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1100_inst_req_1 : boolean;
  signal type_cast_1370_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1100_inst_ack_1 : boolean;
  signal type_cast_1005_inst_ack_1 : boolean;
  signal type_cast_1316_inst_ack_1 : boolean;
  signal type_cast_1104_inst_req_0 : boolean;
  signal type_cast_1104_inst_ack_0 : boolean;
  signal if_stmt_1486_branch_ack_1 : boolean;
  signal type_cast_1104_inst_req_1 : boolean;
  signal type_cast_1104_inst_ack_1 : boolean;
  signal type_cast_1469_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1118_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1118_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1118_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1118_inst_ack_1 : boolean;
  signal type_cast_1316_inst_req_1 : boolean;
  signal type_cast_1122_inst_req_0 : boolean;
  signal type_cast_1122_inst_ack_0 : boolean;
  signal type_cast_1122_inst_req_1 : boolean;
  signal type_cast_1122_inst_ack_1 : boolean;
  signal type_cast_1539_inst_ack_0 : boolean;
  signal type_cast_1469_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1136_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1366_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1136_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1136_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1366_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1136_inst_ack_1 : boolean;
  signal type_cast_1005_inst_req_0 : boolean;
  signal type_cast_1406_inst_ack_1 : boolean;
  signal type_cast_1406_inst_req_1 : boolean;
  signal type_cast_1316_inst_ack_0 : boolean;
  signal if_stmt_1486_branch_req_0 : boolean;
  signal type_cast_1140_inst_req_0 : boolean;
  signal type_cast_1140_inst_ack_0 : boolean;
  signal type_cast_1140_inst_req_1 : boolean;
  signal type_cast_1140_inst_ack_1 : boolean;
  signal type_cast_1515_inst_ack_1 : boolean;
  signal type_cast_1316_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1366_inst_ack_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1312_inst_ack_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1312_inst_req_1 : boolean;
  signal RPIPE_maxpool_input_pipe_1366_inst_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1312_inst_ack_0 : boolean;
  signal ptr_deref_1148_store_0_req_0 : boolean;
  signal RPIPE_maxpool_input_pipe_1312_inst_req_0 : boolean;
  signal ptr_deref_1148_store_0_ack_0 : boolean;
  signal ptr_deref_1148_store_0_req_1 : boolean;
  signal ptr_deref_1148_store_0_ack_1 : boolean;
  signal array_obj_ref_1295_index_offset_ack_1 : boolean;
  signal type_cast_1406_inst_ack_0 : boolean;
  signal array_obj_ref_1295_index_offset_req_1 : boolean;
  signal type_cast_1303_inst_ack_1 : boolean;
  signal type_cast_1303_inst_req_1 : boolean;
  signal type_cast_1462_inst_ack_1 : boolean;
  signal type_cast_1462_inst_req_1 : boolean;
  signal if_stmt_1162_branch_req_0 : boolean;
  signal if_stmt_1162_branch_ack_1 : boolean;
  signal if_stmt_1162_branch_ack_0 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal type_cast_1173_inst_req_1 : boolean;
  signal type_cast_1173_inst_ack_1 : boolean;
  signal phi_stmt_999_req_1 : boolean;
  signal type_cast_1177_inst_req_0 : boolean;
  signal type_cast_1177_inst_ack_0 : boolean;
  signal type_cast_1177_inst_req_1 : boolean;
  signal type_cast_1177_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1852_inst_req_1 : boolean;
  signal if_stmt_1200_branch_req_0 : boolean;
  signal if_stmt_1200_branch_ack_1 : boolean;
  signal if_stmt_1200_branch_ack_0 : boolean;
  signal phi_stmt_1526_req_0 : boolean;
  signal phi_stmt_999_ack_0 : boolean;
  signal type_cast_1221_inst_req_0 : boolean;
  signal type_cast_1221_inst_ack_0 : boolean;
  signal type_cast_1221_inst_req_1 : boolean;
  signal type_cast_1221_inst_ack_1 : boolean;
  signal type_cast_1230_inst_req_0 : boolean;
  signal type_cast_1230_inst_ack_0 : boolean;
  signal type_cast_1230_inst_req_1 : boolean;
  signal type_cast_1230_inst_ack_1 : boolean;
  signal type_cast_1239_inst_req_0 : boolean;
  signal type_cast_1239_inst_ack_0 : boolean;
  signal type_cast_1239_inst_req_1 : boolean;
  signal type_cast_1239_inst_ack_1 : boolean;
  signal type_cast_1273_inst_req_0 : boolean;
  signal type_cast_1273_inst_ack_0 : boolean;
  signal type_cast_1273_inst_req_1 : boolean;
  signal type_cast_1273_inst_ack_1 : boolean;
  signal type_cast_1577_inst_req_0 : boolean;
  signal type_cast_1577_inst_ack_0 : boolean;
  signal type_cast_1577_inst_req_1 : boolean;
  signal type_cast_1577_inst_ack_1 : boolean;
  signal phi_stmt_1519_req_0 : boolean;
  signal type_cast_1522_inst_ack_1 : boolean;
  signal type_cast_1522_inst_req_1 : boolean;
  signal array_obj_ref_1606_index_offset_req_0 : boolean;
  signal array_obj_ref_1606_index_offset_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1852_inst_req_0 : boolean;
  signal array_obj_ref_1606_index_offset_req_1 : boolean;
  signal array_obj_ref_1606_index_offset_ack_1 : boolean;
  signal type_cast_1529_inst_ack_0 : boolean;
  signal phi_stmt_1570_ack_0 : boolean;
  signal addr_of_1607_final_reg_req_0 : boolean;
  signal addr_of_1607_final_reg_ack_0 : boolean;
  signal addr_of_1607_final_reg_req_1 : boolean;
  signal addr_of_1607_final_reg_ack_1 : boolean;
  signal type_cast_1522_inst_ack_0 : boolean;
  signal type_cast_1522_inst_req_0 : boolean;
  signal phi_stmt_1570_req_0 : boolean;
  signal ptr_deref_1610_store_0_req_0 : boolean;
  signal ptr_deref_1610_store_0_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1846_inst_ack_1 : boolean;
  signal ptr_deref_1610_store_0_req_1 : boolean;
  signal ptr_deref_1610_store_0_ack_1 : boolean;
  signal phi_stmt_999_req_0 : boolean;
  signal type_cast_1573_inst_ack_1 : boolean;
  signal call_stmt_1617_call_req_0 : boolean;
  signal call_stmt_1617_call_ack_0 : boolean;
  signal type_cast_1573_inst_req_1 : boolean;
  signal call_stmt_1617_call_req_1 : boolean;
  signal call_stmt_1617_call_ack_1 : boolean;
  signal WPIPE_output_pipe_1618_inst_req_0 : boolean;
  signal WPIPE_output_pipe_1618_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_1618_inst_req_1 : boolean;
  signal WPIPE_output_pipe_1618_inst_ack_1 : boolean;
  signal phi_stmt_1672_ack_0 : boolean;
  signal WPIPE_output_pipe_1621_inst_req_0 : boolean;
  signal WPIPE_output_pipe_1621_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_1621_inst_req_1 : boolean;
  signal WPIPE_output_pipe_1621_inst_ack_1 : boolean;
  signal phi_stmt_1672_req_0 : boolean;
  signal WPIPE_output_pipe_1624_inst_req_0 : boolean;
  signal WPIPE_output_pipe_1624_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_1624_inst_req_1 : boolean;
  signal phi_stmt_1283_ack_0 : boolean;
  signal WPIPE_output_pipe_1624_inst_ack_1 : boolean;
  signal type_cast_1675_inst_ack_1 : boolean;
  signal type_cast_1675_inst_req_1 : boolean;
  signal type_cast_1675_inst_ack_0 : boolean;
  signal type_cast_1529_inst_req_0 : boolean;
  signal type_cast_1573_inst_ack_0 : boolean;
  signal type_cast_1642_inst_req_0 : boolean;
  signal type_cast_1642_inst_ack_0 : boolean;
  signal type_cast_1573_inst_req_0 : boolean;
  signal type_cast_1642_inst_req_1 : boolean;
  signal type_cast_1642_inst_ack_1 : boolean;
  signal type_cast_1663_inst_req_0 : boolean;
  signal phi_stmt_1283_req_1 : boolean;
  signal type_cast_1663_inst_ack_0 : boolean;
  signal type_cast_1663_inst_req_1 : boolean;
  signal type_cast_1289_inst_ack_1 : boolean;
  signal type_cast_1663_inst_ack_1 : boolean;
  signal type_cast_1675_inst_req_0 : boolean;
  signal type_cast_1289_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1685_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1685_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1685_inst_req_1 : boolean;
  signal WPIPE_num_out_pipe_1685_inst_ack_1 : boolean;
  signal WPIPE_num_out_pipe_1688_inst_req_0 : boolean;
  signal type_cast_1289_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1688_inst_ack_0 : boolean;
  signal WPIPE_num_out_pipe_1688_inst_req_1 : boolean;
  signal type_cast_1289_inst_req_0 : boolean;
  signal WPIPE_num_out_pipe_1688_inst_ack_1 : boolean;
  signal call_stmt_1693_call_req_0 : boolean;
  signal call_stmt_1693_call_ack_0 : boolean;
  signal call_stmt_1693_call_req_1 : boolean;
  signal call_stmt_1693_call_ack_1 : boolean;
  signal call_stmt_1697_call_req_0 : boolean;
  signal call_stmt_1697_call_ack_0 : boolean;
  signal call_stmt_1697_call_req_1 : boolean;
  signal call_stmt_1697_call_ack_1 : boolean;
  signal phi_stmt_1466_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1846_inst_req_1 : boolean;
  signal if_stmt_1709_branch_req_0 : boolean;
  signal if_stmt_1709_branch_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1846_inst_ack_0 : boolean;
  signal if_stmt_1709_branch_ack_0 : boolean;
  signal type_cast_1720_inst_req_0 : boolean;
  signal type_cast_1720_inst_ack_0 : boolean;
  signal phi_stmt_1526_ack_0 : boolean;
  signal type_cast_1720_inst_req_1 : boolean;
  signal type_cast_1720_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1723_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_1723_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1849_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_1723_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_1723_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1849_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_1727_inst_req_0 : boolean;
  signal RPIPE_input_done_pipe_1727_inst_ack_0 : boolean;
  signal RPIPE_input_done_pipe_1727_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_1727_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1852_inst_ack_1 : boolean;
  signal phi_stmt_1466_req_1 : boolean;
  signal call_stmt_1731_call_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1858_inst_req_0 : boolean;
  signal call_stmt_1731_call_ack_0 : boolean;
  signal phi_stmt_1519_ack_0 : boolean;
  signal call_stmt_1731_call_req_1 : boolean;
  signal call_stmt_1731_call_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1843_inst_ack_1 : boolean;
  signal phi_stmt_1283_req_0 : boolean;
  signal type_cast_1735_inst_req_0 : boolean;
  signal type_cast_1735_inst_ack_0 : boolean;
  signal phi_stmt_1526_req_1 : boolean;
  signal type_cast_1735_inst_req_1 : boolean;
  signal type_cast_1735_inst_ack_1 : boolean;
  signal type_cast_1744_inst_req_0 : boolean;
  signal type_cast_1744_inst_ack_0 : boolean;
  signal phi_stmt_1672_req_1 : boolean;
  signal type_cast_1744_inst_req_1 : boolean;
  signal type_cast_1744_inst_ack_1 : boolean;
  signal phi_stmt_1466_req_0 : boolean;
  signal type_cast_1748_inst_req_0 : boolean;
  signal type_cast_1748_inst_ack_0 : boolean;
  signal type_cast_1748_inst_req_1 : boolean;
  signal type_cast_1748_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1843_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1849_inst_ack_0 : boolean;
  signal type_cast_1469_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_ack_1 : boolean;
  signal call_stmt_1761_call_req_0 : boolean;
  signal call_stmt_1761_call_ack_0 : boolean;
  signal phi_stmt_1519_req_1 : boolean;
  signal call_stmt_1761_call_req_1 : boolean;
  signal call_stmt_1761_call_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1849_inst_req_0 : boolean;
  signal type_cast_1469_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1855_inst_req_1 : boolean;
  signal type_cast_1765_inst_req_0 : boolean;
  signal type_cast_1765_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1846_inst_req_0 : boolean;
  signal type_cast_1765_inst_req_1 : boolean;
  signal type_cast_1765_inst_ack_1 : boolean;
  signal type_cast_1775_inst_req_0 : boolean;
  signal type_cast_1775_inst_ack_0 : boolean;
  signal type_cast_1775_inst_req_1 : boolean;
  signal type_cast_1775_inst_ack_1 : boolean;
  signal type_cast_1785_inst_req_0 : boolean;
  signal type_cast_1785_inst_ack_0 : boolean;
  signal type_cast_1785_inst_req_1 : boolean;
  signal type_cast_1785_inst_ack_1 : boolean;
  signal type_cast_1795_inst_req_0 : boolean;
  signal type_cast_1795_inst_ack_0 : boolean;
  signal type_cast_1795_inst_req_1 : boolean;
  signal type_cast_1795_inst_ack_1 : boolean;
  signal type_cast_1805_inst_req_0 : boolean;
  signal type_cast_1805_inst_ack_0 : boolean;
  signal type_cast_1805_inst_req_1 : boolean;
  signal type_cast_1805_inst_ack_1 : boolean;
  signal type_cast_1815_inst_req_0 : boolean;
  signal type_cast_1815_inst_ack_0 : boolean;
  signal type_cast_1815_inst_req_1 : boolean;
  signal type_cast_1815_inst_ack_1 : boolean;
  signal type_cast_1825_inst_req_0 : boolean;
  signal type_cast_1825_inst_ack_0 : boolean;
  signal type_cast_1825_inst_req_1 : boolean;
  signal type_cast_1825_inst_ack_1 : boolean;
  signal type_cast_1835_inst_req_0 : boolean;
  signal type_cast_1835_inst_ack_0 : boolean;
  signal type_cast_1835_inst_req_1 : boolean;
  signal type_cast_1835_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1837_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1840_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1840_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1840_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1840_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_1843_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_1843_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolution3D_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolution3D_CP_2151_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolution3D_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_2151_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolution3D_CP_2151_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolution3D_CP_2151_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolution3D_CP_2151: Block -- control-path 
    signal convolution3D_CP_2151_elements: BooleanArray(326 downto 0);
    -- 
  begin -- 
    convolution3D_CP_2151_elements(0) <= convolution3D_CP_2151_start;
    convolution3D_CP_2151_symbol <= convolution3D_CP_2151_elements(282);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	40 
    -- CP-element group 0: 	44 
    -- CP-element group 0: 	48 
    -- CP-element group 0: 	28 
    -- CP-element group 0: 	32 
    -- CP-element group 0: 	36 
    -- CP-element group 0: 	16 
    -- CP-element group 0: 	20 
    -- CP-element group 0: 	24 
    -- CP-element group 0: 	64 
    -- CP-element group 0: 	67 
    -- CP-element group 0: 	70 
    -- CP-element group 0: 	52 
    -- CP-element group 0: 	56 
    -- CP-element group 0: 	60 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	8 
    -- CP-element group 0: 	12 
    -- CP-element group 0:  members (62) 
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Update/cr
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_720/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/branch_block_stmt_720__entry__
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944__entry__
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_update_start_
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Update/cr
      -- 
    cr_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_814_inst_req_1); -- 
    rr_2249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => RPIPE_maxpool_input_pipe_722_inst_req_0); -- 
    cr_2268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_726_inst_req_1); -- 
    cr_2324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_751_inst_req_1); -- 
    cr_2520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_839_inst_req_1); -- 
    cr_2492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_826_inst_req_1); -- 
    cr_2548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_851_inst_req_1); -- 
    cr_2436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_801_inst_req_1); -- 
    cr_2352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_764_inst_req_1); -- 
    cr_2576_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2576_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_864_inst_req_1); -- 
    cr_2632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_889_inst_req_1); -- 
    cr_2380_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2380_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_776_inst_req_1); -- 
    cr_2296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_739_inst_req_1); -- 
    cr_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_876_inst_req_1); -- 
    cr_2408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_789_inst_req_1); -- 
    cr_2660_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2660_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_901_inst_req_1); -- 
    cr_2688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_914_inst_req_1); -- 
    cr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2702_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_923_inst_req_1); -- 
    cr_2716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(0), ack => type_cast_927_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_update_start_
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Sample/ra
      -- 
    ra_2250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_722_inst_ack_0, ack => convolution3D_CP_2151_elements(1)); -- 
    cr_2254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(1), ack => RPIPE_maxpool_input_pipe_722_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_722_update_completed_
      -- 
    ca_2255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_722_inst_ack_1, ack => convolution3D_CP_2151_elements(2)); -- 
    rr_2263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(2), ack => type_cast_726_inst_req_0); -- 
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(2), ack => RPIPE_maxpool_input_pipe_735_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_sample_completed_
      -- 
    ra_2264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_726_inst_ack_0, ack => convolution3D_CP_2151_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	71 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_726_update_completed_
      -- 
    ca_2269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_726_inst_ack_1, ack => convolution3D_CP_2151_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_update_start_
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Update/cr
      -- CP-element group 5: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Update/$entry
      -- 
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_735_inst_ack_0, ack => convolution3D_CP_2151_elements(5)); -- 
    cr_2282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(5), ack => RPIPE_maxpool_input_pipe_735_inst_req_1); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Update/ca
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_735_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Sample/rr
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_sample_start_
      -- 
    ca_2283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_735_inst_ack_1, ack => convolution3D_CP_2151_elements(6)); -- 
    rr_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(6), ack => type_cast_739_inst_req_0); -- 
    rr_2305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(6), ack => RPIPE_maxpool_input_pipe_747_inst_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_sample_completed_
      -- 
    ra_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_0, ack => convolution3D_CP_2151_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	0 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	71 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_739_Update/$exit
      -- 
    ca_2297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_739_inst_ack_1, ack => convolution3D_CP_2151_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Update/cr
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_update_start_
      -- CP-element group 9: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_sample_completed_
      -- 
    ra_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_747_inst_ack_0, ack => convolution3D_CP_2151_elements(9)); -- 
    cr_2310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(9), ack => RPIPE_maxpool_input_pipe_747_inst_req_1); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Update/ca
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_747_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Sample/$entry
      -- 
    ca_2311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_747_inst_ack_1, ack => convolution3D_CP_2151_elements(10)); -- 
    rr_2319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(10), ack => type_cast_751_inst_req_0); -- 
    rr_2333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(10), ack => RPIPE_maxpool_input_pipe_760_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Sample/$exit
      -- 
    ra_2320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => convolution3D_CP_2151_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	0 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	65 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_751_Update/$exit
      -- 
    ca_2325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_1, ack => convolution3D_CP_2151_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_update_start_
      -- CP-element group 13: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_sample_completed_
      -- 
    ra_2334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_760_inst_ack_0, ack => convolution3D_CP_2151_elements(13)); -- 
    cr_2338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(13), ack => RPIPE_maxpool_input_pipe_760_inst_req_1); -- 
    -- CP-element group 14:  fork  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	17 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_760_update_completed_
      -- 
    ca_2339_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_760_inst_ack_1, ack => convolution3D_CP_2151_elements(14)); -- 
    rr_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(14), ack => type_cast_764_inst_req_0); -- 
    rr_2361_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2361_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(14), ack => RPIPE_maxpool_input_pipe_772_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Sample/ra
      -- 
    ra_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_0, ack => convolution3D_CP_2151_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	0 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	65 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_764_Update/$exit
      -- 
    ca_2353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_764_inst_ack_1, ack => convolution3D_CP_2151_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_update_start_
      -- CP-element group 17: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_sample_completed_
      -- 
    ra_2362_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_772_inst_ack_0, ack => convolution3D_CP_2151_elements(17)); -- 
    cr_2366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(17), ack => RPIPE_maxpool_input_pipe_772_inst_req_1); -- 
    -- CP-element group 18:  fork  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_772_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Sample/rr
      -- CP-element group 18: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Sample/$entry
      -- 
    ca_2367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_772_inst_ack_1, ack => convolution3D_CP_2151_elements(18)); -- 
    rr_2375_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2375_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(18), ack => type_cast_776_inst_req_0); -- 
    rr_2389_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2389_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(18), ack => RPIPE_maxpool_input_pipe_785_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Sample/$exit
      -- 
    ra_2376_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_0, ack => convolution3D_CP_2151_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	0 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	68 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_776_update_completed_
      -- 
    ca_2381_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_776_inst_ack_1, ack => convolution3D_CP_2151_elements(20)); -- 
    -- CP-element group 21:  transition  input  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (6) 
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Update/cr
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_update_start_
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Update/$entry
      -- 
    ra_2390_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_785_inst_ack_0, ack => convolution3D_CP_2151_elements(21)); -- 
    cr_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(21), ack => RPIPE_maxpool_input_pipe_785_inst_req_1); -- 
    -- CP-element group 22:  fork  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	25 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Sample/rr
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_785_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_sample_start_
      -- 
    ca_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_785_inst_ack_1, ack => convolution3D_CP_2151_elements(22)); -- 
    rr_2403_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2403_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(22), ack => type_cast_789_inst_req_0); -- 
    rr_2417_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2417_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(22), ack => RPIPE_maxpool_input_pipe_797_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Sample/ra
      -- CP-element group 23: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_sample_completed_
      -- 
    ra_2404_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_789_inst_ack_0, ack => convolution3D_CP_2151_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	0 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	68 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_789_Update/$exit
      -- 
    ca_2409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_789_inst_ack_1, ack => convolution3D_CP_2151_elements(24)); -- 
    -- CP-element group 25:  transition  input  output  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	22 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	26 
    -- CP-element group 25:  members (6) 
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Update/cr
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_update_start_
      -- CP-element group 25: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_sample_completed_
      -- 
    ra_2418_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_797_inst_ack_0, ack => convolution3D_CP_2151_elements(25)); -- 
    cr_2422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(25), ack => RPIPE_maxpool_input_pipe_797_inst_req_1); -- 
    -- CP-element group 26:  fork  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	25 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Sample/rr
      -- CP-element group 26: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_797_update_completed_
      -- 
    ca_2423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_797_inst_ack_1, ack => convolution3D_CP_2151_elements(26)); -- 
    rr_2431_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2431_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(26), ack => type_cast_801_inst_req_0); -- 
    rr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(26), ack => RPIPE_maxpool_input_pipe_810_inst_req_0); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_sample_completed_
      -- 
    ra_2432_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_0, ack => convolution3D_CP_2151_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	0 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	71 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_801_Update/$exit
      -- 
    ca_2437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_801_inst_ack_1, ack => convolution3D_CP_2151_elements(28)); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	26 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_update_start_
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Sample/ra
      -- 
    ra_2446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_0, ack => convolution3D_CP_2151_elements(29)); -- 
    cr_2450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(29), ack => RPIPE_maxpool_input_pipe_810_inst_req_1); -- 
    -- CP-element group 30:  fork  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Update/ca
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_810_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Sample/rr
      -- CP-element group 30: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Sample/$entry
      -- 
    ca_2451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_810_inst_ack_1, ack => convolution3D_CP_2151_elements(30)); -- 
    rr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(30), ack => type_cast_814_inst_req_0); -- 
    rr_2473_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2473_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(30), ack => RPIPE_maxpool_input_pipe_822_inst_req_0); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Sample/ra
      -- CP-element group 31: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Sample/$exit
      -- 
    ra_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_0, ack => convolution3D_CP_2151_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	0 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	71 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_Update/ca
      -- CP-element group 32: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_814_update_completed_
      -- 
    ca_2465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_814_inst_ack_1, ack => convolution3D_CP_2151_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	30 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Update/cr
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Sample/ra
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Sample/$exit
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_update_start_
      -- CP-element group 33: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_sample_completed_
      -- 
    ra_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_822_inst_ack_0, ack => convolution3D_CP_2151_elements(33)); -- 
    cr_2478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(33), ack => RPIPE_maxpool_input_pipe_822_inst_req_1); -- 
    -- CP-element group 34:  fork  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	37 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (9) 
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Sample/rr
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Update/ca
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_822_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Sample/$entry
      -- 
    ca_2479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_822_inst_ack_1, ack => convolution3D_CP_2151_elements(34)); -- 
    rr_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(34), ack => type_cast_826_inst_req_0); -- 
    rr_2501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(34), ack => RPIPE_maxpool_input_pipe_835_inst_req_0); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_sample_completed_
      -- 
    ra_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_0, ack => convolution3D_CP_2151_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	0 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	71 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_826_Update/ca
      -- 
    ca_2493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_826_inst_ack_1, ack => convolution3D_CP_2151_elements(36)); -- 
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	34 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Update/cr
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_update_start_
      -- CP-element group 37: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Sample/$exit
      -- 
    ra_2502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_835_inst_ack_0, ack => convolution3D_CP_2151_elements(37)); -- 
    cr_2506_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2506_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(37), ack => RPIPE_maxpool_input_pipe_835_inst_req_1); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: 	41 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_835_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Sample/rr
      -- 
    ca_2507_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_835_inst_ack_1, ack => convolution3D_CP_2151_elements(38)); -- 
    rr_2515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(38), ack => type_cast_839_inst_req_0); -- 
    rr_2529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(38), ack => RPIPE_maxpool_input_pipe_847_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Sample/ra
      -- CP-element group 39: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Sample/$exit
      -- 
    ra_2516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_0, ack => convolution3D_CP_2151_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	0 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	71 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_839_update_completed_
      -- 
    ca_2521_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_839_inst_ack_1, ack => convolution3D_CP_2151_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	38 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (6) 
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Sample/ra
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_update_start_
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Update/cr
      -- 
    ra_2530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_0, ack => convolution3D_CP_2151_elements(41)); -- 
    cr_2534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(41), ack => RPIPE_maxpool_input_pipe_847_inst_req_1); -- 
    -- CP-element group 42:  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: 	45 
    -- CP-element group 42:  members (9) 
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Sample/rr
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_847_Update/ca
      -- 
    ca_2535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_847_inst_ack_1, ack => convolution3D_CP_2151_elements(42)); -- 
    rr_2543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(42), ack => type_cast_851_inst_req_0); -- 
    rr_2557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(42), ack => RPIPE_maxpool_input_pipe_860_inst_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Sample/ra
      -- CP-element group 43: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_sample_completed_
      -- 
    ra_2544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_0, ack => convolution3D_CP_2151_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	0 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	71 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Update/ca
      -- CP-element group 44: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_851_Update/$exit
      -- 
    ca_2549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_851_inst_ack_1, ack => convolution3D_CP_2151_elements(44)); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	42 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Update/cr
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_update_start_
      -- CP-element group 45: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Sample/$exit
      -- 
    ra_2558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_860_inst_ack_0, ack => convolution3D_CP_2151_elements(45)); -- 
    cr_2562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(45), ack => RPIPE_maxpool_input_pipe_860_inst_req_1); -- 
    -- CP-element group 46:  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46: 	49 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_860_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_sample_start_
      -- 
    ca_2563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_860_inst_ack_1, ack => convolution3D_CP_2151_elements(46)); -- 
    rr_2571_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2571_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(46), ack => type_cast_864_inst_req_0); -- 
    rr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2585_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(46), ack => RPIPE_maxpool_input_pipe_872_inst_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Sample/ra
      -- CP-element group 47: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Sample/$exit
      -- 
    ra_2572_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_0, ack => convolution3D_CP_2151_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	0 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	71 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_864_Update/ca
      -- 
    ca_2577_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_864_inst_ack_1, ack => convolution3D_CP_2151_elements(48)); -- 
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	46 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Update/cr
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Sample/ra
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_update_start_
      -- 
    ra_2586_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_872_inst_ack_0, ack => convolution3D_CP_2151_elements(49)); -- 
    cr_2590_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2590_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(49), ack => RPIPE_maxpool_input_pipe_872_inst_req_1); -- 
    -- CP-element group 50:  fork  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	53 
    -- CP-element group 50:  members (9) 
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_872_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Sample/rr
      -- 
    ca_2591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_872_inst_ack_1, ack => convolution3D_CP_2151_elements(50)); -- 
    rr_2599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(50), ack => type_cast_876_inst_req_0); -- 
    rr_2613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(50), ack => RPIPE_maxpool_input_pipe_885_inst_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Sample/ra
      -- 
    ra_2600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_876_inst_ack_0, ack => convolution3D_CP_2151_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	0 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	71 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_876_Update/$exit
      -- 
    ca_2605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_876_inst_ack_1, ack => convolution3D_CP_2151_elements(52)); -- 
    -- CP-element group 53:  transition  input  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	50 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (6) 
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Update/$entry
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Update/cr
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_update_start_
      -- CP-element group 53: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Sample/ra
      -- 
    ra_2614_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_885_inst_ack_0, ack => convolution3D_CP_2151_elements(53)); -- 
    cr_2618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(53), ack => RPIPE_maxpool_input_pipe_885_inst_req_1); -- 
    -- CP-element group 54:  fork  transition  input  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: 	57 
    -- CP-element group 54:  members (9) 
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_885_update_completed_
      -- 
    ca_2619_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_885_inst_ack_1, ack => convolution3D_CP_2151_elements(54)); -- 
    rr_2627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(54), ack => type_cast_889_inst_req_0); -- 
    rr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(54), ack => RPIPE_maxpool_input_pipe_897_inst_req_0); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Sample/ra
      -- CP-element group 55: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_sample_completed_
      -- 
    ra_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_889_inst_ack_0, ack => convolution3D_CP_2151_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	0 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	71 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_Update/ca
      -- CP-element group 56: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_889_update_completed_
      -- 
    ca_2633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_889_inst_ack_1, ack => convolution3D_CP_2151_elements(56)); -- 
    -- CP-element group 57:  transition  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	54 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (6) 
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_update_start_
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Sample/ra
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Update/cr
      -- 
    ra_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_897_inst_ack_0, ack => convolution3D_CP_2151_elements(57)); -- 
    cr_2646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(57), ack => RPIPE_maxpool_input_pipe_897_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	61 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (9) 
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_897_Update/ca
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Sample/rr
      -- 
    ca_2647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_897_inst_ack_1, ack => convolution3D_CP_2151_elements(58)); -- 
    rr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(58), ack => RPIPE_maxpool_input_pipe_910_inst_req_0); -- 
    rr_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(58), ack => type_cast_901_inst_req_0); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Sample/ra
      -- 
    ra_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_0, ack => convolution3D_CP_2151_elements(59)); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	0 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	71 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_901_Update/ca
      -- 
    ca_2661_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_901_inst_ack_1, ack => convolution3D_CP_2151_elements(60)); -- 
    -- CP-element group 61:  transition  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	58 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_update_start_
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Update/cr
      -- 
    ra_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_910_inst_ack_0, ack => convolution3D_CP_2151_elements(61)); -- 
    cr_2674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(61), ack => RPIPE_maxpool_input_pipe_910_inst_req_1); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/RPIPE_maxpool_input_pipe_910_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Sample/rr
      -- 
    ca_2675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_910_inst_ack_1, ack => convolution3D_CP_2151_elements(62)); -- 
    rr_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(62), ack => type_cast_914_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Sample/ra
      -- 
    ra_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_0, ack => convolution3D_CP_2151_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	0 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	71 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_914_Update/ca
      -- 
    ca_2689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_1, ack => convolution3D_CP_2151_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	16 
    -- CP-element group 65: 	12 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Sample/rr
      -- 
    rr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(65), ack => type_cast_923_inst_req_0); -- 
    convolution3D_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(16) & convolution3D_CP_2151_elements(12);
      gj_convolution3D_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  transition  input  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Sample/ra
      -- 
    ra_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => convolution3D_CP_2151_elements(66)); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	0 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	71 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_923_Update/ca
      -- 
    ca_2703_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_1, ack => convolution3D_CP_2151_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	20 
    -- CP-element group 68: 	24 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Sample/rr
      -- 
    rr_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(68), ack => type_cast_927_inst_req_0); -- 
    convolution3D_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(20) & convolution3D_CP_2151_elements(24);
      gj_convolution3D_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Sample/ra
      -- 
    ra_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_0, ack => convolution3D_CP_2151_elements(69)); -- 
    -- CP-element group 70:  transition  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	0 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/type_cast_927_Update/ca
      -- 
    ca_2717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_927_inst_ack_1, ack => convolution3D_CP_2151_elements(70)); -- 
    -- CP-element group 71:  branch  join  transition  place  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	40 
    -- CP-element group 71: 	44 
    -- CP-element group 71: 	48 
    -- CP-element group 71: 	28 
    -- CP-element group 71: 	32 
    -- CP-element group 71: 	36 
    -- CP-element group 71: 	64 
    -- CP-element group 71: 	67 
    -- CP-element group 71: 	70 
    -- CP-element group 71: 	52 
    -- CP-element group 71: 	56 
    -- CP-element group 71: 	60 
    -- CP-element group 71: 	4 
    -- CP-element group 71: 	8 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (10) 
      -- CP-element group 71: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944/$exit
      -- CP-element group 71: 	 branch_block_stmt_720/assign_stmt_723_to_assign_stmt_944__exit__
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945__entry__
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_dead_link/$entry
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_eval_test/$entry
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_eval_test/$exit
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_eval_test/branch_req
      -- CP-element group 71: 	 branch_block_stmt_720/R_cmp343_946_place
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_if_link/$entry
      -- CP-element group 71: 	 branch_block_stmt_720/if_stmt_945_else_link/$entry
      -- 
    branch_req_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(71), ack => if_stmt_945_branch_req_0); -- 
    convolution3D_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 33) := "convolution3D_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(40) & convolution3D_CP_2151_elements(44) & convolution3D_CP_2151_elements(48) & convolution3D_CP_2151_elements(28) & convolution3D_CP_2151_elements(32) & convolution3D_CP_2151_elements(36) & convolution3D_CP_2151_elements(64) & convolution3D_CP_2151_elements(67) & convolution3D_CP_2151_elements(70) & convolution3D_CP_2151_elements(52) & convolution3D_CP_2151_elements(56) & convolution3D_CP_2151_elements(60) & convolution3D_CP_2151_elements(4) & convolution3D_CP_2151_elements(8);
      gj_convolution3D_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: 	75 
    -- CP-element group 72:  members (18) 
      -- CP-element group 72: 	 branch_block_stmt_720/merge_stmt_951__exit__
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996__entry__
      -- CP-element group 72: 	 branch_block_stmt_720/if_stmt_945_if_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_720/if_stmt_945_if_link/if_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_720/entry_bbx_xnph345
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/$entry
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_update_start_
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Update/cr
      -- CP-element group 72: 	 branch_block_stmt_720/merge_stmt_951_PhiAck/dummy
      -- CP-element group 72: 	 branch_block_stmt_720/merge_stmt_951_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_720/merge_stmt_951_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_720/entry_bbx_xnph345_PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_720/entry_bbx_xnph345_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_720/merge_stmt_951_PhiReqMerge
      -- 
    if_choice_transition_2730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_945_branch_ack_1, ack => convolution3D_CP_2151_elements(72)); -- 
    rr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(72), ack => type_cast_982_inst_req_0); -- 
    cr_2752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(72), ack => type_cast_982_inst_req_1); -- 
    -- CP-element group 73:  transition  place  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	289 
    -- CP-element group 73:  members (5) 
      -- CP-element group 73: 	 branch_block_stmt_720/if_stmt_945_else_link/$exit
      -- CP-element group 73: 	 branch_block_stmt_720/if_stmt_945_else_link/else_choice_transition
      -- CP-element group 73: 	 branch_block_stmt_720/entry_forx_xend
      -- CP-element group 73: 	 branch_block_stmt_720/entry_forx_xend_PhiReq/$exit
      -- CP-element group 73: 	 branch_block_stmt_720/entry_forx_xend_PhiReq/$entry
      -- 
    else_choice_transition_2734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_945_branch_ack_0, ack => convolution3D_CP_2151_elements(73)); -- 
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Sample/ra
      -- 
    ra_2748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_982_inst_ack_0, ack => convolution3D_CP_2151_elements(74)); -- 
    -- CP-element group 75:  transition  place  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	72 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	283 
    -- CP-element group 75:  members (9) 
      -- CP-element group 75: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996__exit__
      -- CP-element group 75: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody
      -- CP-element group 75: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/$exit
      -- CP-element group 75: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_720/assign_stmt_956_to_assign_stmt_996/type_cast_982_Update/ca
      -- CP-element group 75: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/$entry
      -- CP-element group 75: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/$entry
      -- CP-element group 75: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/$entry
      -- 
    ca_2753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_982_inst_ack_1, ack => convolution3D_CP_2151_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	288 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	115 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_sample_complete
      -- CP-element group 76: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Sample/ack
      -- 
    ack_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1011_index_offset_ack_0, ack => convolution3D_CP_2151_elements(76)); -- 
    -- CP-element group 77:  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	288 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (11) 
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_root_address_calculated
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_offset_calculated
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Update/ack
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_base_plus_offset/$entry
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_base_plus_offset/$exit
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_base_plus_offset/sum_rename_req
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_base_plus_offset/sum_rename_ack
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_request/$entry
      -- CP-element group 77: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_request/req
      -- 
    ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1011_index_offset_ack_1, ack => convolution3D_CP_2151_elements(77)); -- 
    req_2796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(77), ack => addr_of_1012_final_reg_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_request/$exit
      -- CP-element group 78: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_request/ack
      -- 
    ack_2797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1012_final_reg_ack_0, ack => convolution3D_CP_2151_elements(78)); -- 
    -- CP-element group 79:  fork  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	288 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	112 
    -- CP-element group 79:  members (19) 
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_complete/$exit
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_complete/ack
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_address_calculated
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_word_address_calculated
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_root_address_calculated
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_address_resized
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_addr_resize/$entry
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_addr_resize/$exit
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_addr_resize/base_resize_req
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_addr_resize/base_resize_ack
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_plus_offset/$entry
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_plus_offset/$exit
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_plus_offset/sum_rename_req
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_base_plus_offset/sum_rename_ack
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_word_addrgen/$entry
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_word_addrgen/$exit
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_word_addrgen/root_register_req
      -- CP-element group 79: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_word_addrgen/root_register_ack
      -- 
    ack_2802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1012_final_reg_ack_1, ack => convolution3D_CP_2151_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	288 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_update_start_
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Sample/ra
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Update/$entry
      -- CP-element group 80: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Update/cr
      -- 
    ra_2811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1015_inst_ack_0, ack => convolution3D_CP_2151_elements(80)); -- 
    cr_2815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(80), ack => RPIPE_maxpool_input_pipe_1015_inst_req_1); -- 
    -- CP-element group 81:  fork  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	84 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (9) 
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Update/ca
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Sample/rr
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_sample_start_
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Sample/$entry
      -- CP-element group 81: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Sample/rr
      -- 
    ca_2816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1015_inst_ack_1, ack => convolution3D_CP_2151_elements(81)); -- 
    rr_2838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(81), ack => RPIPE_maxpool_input_pipe_1028_inst_req_0); -- 
    rr_2824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(81), ack => type_cast_1019_inst_req_0); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Sample/ra
      -- 
    ra_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_0, ack => convolution3D_CP_2151_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	288 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	112 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Update/ca
      -- 
    ca_2830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1019_inst_ack_1, ack => convolution3D_CP_2151_elements(83)); -- 
    -- CP-element group 84:  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	81 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (6) 
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_update_start_
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Sample/ra
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Update/cr
      -- 
    ra_2839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1028_inst_ack_0, ack => convolution3D_CP_2151_elements(84)); -- 
    cr_2843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(84), ack => RPIPE_maxpool_input_pipe_1028_inst_req_1); -- 
    -- CP-element group 85:  fork  transition  input  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	88 
    -- CP-element group 85:  members (9) 
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1028_Update/ca
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Sample/rr
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_sample_start_
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Sample/$entry
      -- CP-element group 85: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Sample/rr
      -- 
    ca_2844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1028_inst_ack_1, ack => convolution3D_CP_2151_elements(85)); -- 
    rr_2852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(85), ack => type_cast_1032_inst_req_0); -- 
    rr_2866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(85), ack => RPIPE_maxpool_input_pipe_1046_inst_req_0); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Sample/ra
      -- 
    ra_2853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1032_inst_ack_0, ack => convolution3D_CP_2151_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	288 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	112 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Update/ca
      -- 
    ca_2858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1032_inst_ack_1, ack => convolution3D_CP_2151_elements(87)); -- 
    -- CP-element group 88:  transition  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	85 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (6) 
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_update_start_
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Sample/ra
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Update/cr
      -- 
    ra_2867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1046_inst_ack_0, ack => convolution3D_CP_2151_elements(88)); -- 
    cr_2871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(88), ack => RPIPE_maxpool_input_pipe_1046_inst_req_1); -- 
    -- CP-element group 89:  fork  transition  input  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	92 
    -- CP-element group 89:  members (9) 
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1046_Update/ca
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Sample/rr
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Sample/$entry
      -- CP-element group 89: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Sample/rr
      -- 
    ca_2872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1046_inst_ack_1, ack => convolution3D_CP_2151_elements(89)); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(89), ack => type_cast_1050_inst_req_0); -- 
    rr_2894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(89), ack => RPIPE_maxpool_input_pipe_1064_inst_req_0); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Sample/ra
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_0, ack => convolution3D_CP_2151_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	288 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	112 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Update/ca
      -- 
    ca_2886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1050_inst_ack_1, ack => convolution3D_CP_2151_elements(91)); -- 
    -- CP-element group 92:  transition  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	89 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (6) 
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_update_start_
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Update/cr
      -- 
    ra_2895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1064_inst_ack_0, ack => convolution3D_CP_2151_elements(92)); -- 
    cr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(92), ack => RPIPE_maxpool_input_pipe_1064_inst_req_1); -- 
    -- CP-element group 93:  fork  transition  input  output  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93: 	96 
    -- CP-element group 93:  members (9) 
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1064_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Sample/rr
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Sample/$entry
      -- CP-element group 93: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Sample/rr
      -- 
    ca_2900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1064_inst_ack_1, ack => convolution3D_CP_2151_elements(93)); -- 
    rr_2908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(93), ack => type_cast_1068_inst_req_0); -- 
    rr_2922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(93), ack => RPIPE_maxpool_input_pipe_1082_inst_req_0); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Sample/ra
      -- 
    ra_2909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1068_inst_ack_0, ack => convolution3D_CP_2151_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	288 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	112 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Update/ca
      -- 
    ca_2914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1068_inst_ack_1, ack => convolution3D_CP_2151_elements(95)); -- 
    -- CP-element group 96:  transition  input  output  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	93 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (6) 
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_sample_completed_
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_update_start_
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Sample/$exit
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Sample/ra
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Update/cr
      -- 
    ra_2923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1082_inst_ack_0, ack => convolution3D_CP_2151_elements(96)); -- 
    cr_2927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(96), ack => RPIPE_maxpool_input_pipe_1082_inst_req_1); -- 
    -- CP-element group 97:  fork  transition  input  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97: 	100 
    -- CP-element group 97:  members (9) 
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_update_completed_
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Update/$exit
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1082_Update/ca
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Sample/rr
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Sample/$entry
      -- CP-element group 97: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Sample/rr
      -- 
    ca_2928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1082_inst_ack_1, ack => convolution3D_CP_2151_elements(97)); -- 
    rr_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(97), ack => type_cast_1086_inst_req_0); -- 
    rr_2950_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2950_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(97), ack => RPIPE_maxpool_input_pipe_1100_inst_req_0); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Sample/ra
      -- 
    ra_2937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1086_inst_ack_0, ack => convolution3D_CP_2151_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	288 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	112 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Update/ca
      -- 
    ca_2942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1086_inst_ack_1, ack => convolution3D_CP_2151_elements(99)); -- 
    -- CP-element group 100:  transition  input  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	97 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_sample_completed_
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_update_start_
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Sample/ra
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Update/cr
      -- 
    ra_2951_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1100_inst_ack_0, ack => convolution3D_CP_2151_elements(100)); -- 
    cr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(100), ack => RPIPE_maxpool_input_pipe_1100_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	102 
    -- CP-element group 101: 	104 
    -- CP-element group 101:  members (9) 
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Update/$exit
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1100_Update/ca
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Sample/rr
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Sample/rr
      -- 
    ca_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1100_inst_ack_1, ack => convolution3D_CP_2151_elements(101)); -- 
    rr_2964_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2964_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(101), ack => type_cast_1104_inst_req_0); -- 
    rr_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(101), ack => RPIPE_maxpool_input_pipe_1118_inst_req_0); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	101 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_sample_completed_
      -- CP-element group 102: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Sample/ra
      -- 
    ra_2965_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_0, ack => convolution3D_CP_2151_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	288 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	112 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_update_completed_
      -- CP-element group 103: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Update/ca
      -- 
    ca_2970_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1104_inst_ack_1, ack => convolution3D_CP_2151_elements(103)); -- 
    -- CP-element group 104:  transition  input  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	101 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (6) 
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_update_start_
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Update/cr
      -- 
    ra_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1118_inst_ack_0, ack => convolution3D_CP_2151_elements(104)); -- 
    cr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(104), ack => RPIPE_maxpool_input_pipe_1118_inst_req_1); -- 
    -- CP-element group 105:  fork  transition  input  output  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105:  members (9) 
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1118_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Sample/rr
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Sample/$entry
      -- CP-element group 105: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Sample/rr
      -- 
    ca_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1118_inst_ack_1, ack => convolution3D_CP_2151_elements(105)); -- 
    rr_2992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(105), ack => type_cast_1122_inst_req_0); -- 
    rr_3006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(105), ack => RPIPE_maxpool_input_pipe_1136_inst_req_0); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Sample/ra
      -- 
    ra_2993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1122_inst_ack_0, ack => convolution3D_CP_2151_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	288 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	112 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Update/ca
      -- 
    ca_2998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1122_inst_ack_1, ack => convolution3D_CP_2151_elements(107)); -- 
    -- CP-element group 108:  transition  input  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	105 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (6) 
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_update_start_
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Sample/$exit
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Sample/ra
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Update/cr
      -- 
    ra_3007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1136_inst_ack_0, ack => convolution3D_CP_2151_elements(108)); -- 
    cr_3011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(108), ack => RPIPE_maxpool_input_pipe_1136_inst_req_1); -- 
    -- CP-element group 109:  transition  input  output  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109:  members (6) 
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_update_completed_
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1136_Update/ca
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Sample/$entry
      -- CP-element group 109: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Sample/rr
      -- 
    ca_3012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1136_inst_ack_1, ack => convolution3D_CP_2151_elements(109)); -- 
    rr_3020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(109), ack => type_cast_1140_inst_req_0); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Sample/ra
      -- 
    ra_3021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_0, ack => convolution3D_CP_2151_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	288 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Update/ca
      -- 
    ca_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1140_inst_ack_1, ack => convolution3D_CP_2151_elements(111)); -- 
    -- CP-element group 112:  join  transition  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	83 
    -- CP-element group 112: 	87 
    -- CP-element group 112: 	91 
    -- CP-element group 112: 	95 
    -- CP-element group 112: 	99 
    -- CP-element group 112: 	103 
    -- CP-element group 112: 	107 
    -- CP-element group 112: 	111 
    -- CP-element group 112: 	79 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (9) 
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/ptr_deref_1148_Split/$entry
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/ptr_deref_1148_Split/$exit
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/ptr_deref_1148_Split/split_req
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/ptr_deref_1148_Split/split_ack
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/$entry
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/word_0/$entry
      -- CP-element group 112: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/word_0/rr
      -- 
    rr_3064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(112), ack => ptr_deref_1148_store_0_req_0); -- 
    convolution3D_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(83) & convolution3D_CP_2151_elements(87) & convolution3D_CP_2151_elements(91) & convolution3D_CP_2151_elements(95) & convolution3D_CP_2151_elements(99) & convolution3D_CP_2151_elements(103) & convolution3D_CP_2151_elements(107) & convolution3D_CP_2151_elements(111) & convolution3D_CP_2151_elements(79);
      gj_convolution3D_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (5) 
      -- CP-element group 113: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/$exit
      -- CP-element group 113: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Sample/word_access_start/word_0/ra
      -- 
    ra_3065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1148_store_0_ack_0, ack => convolution3D_CP_2151_elements(113)); -- 
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	288 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (5) 
      -- CP-element group 114: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/$exit
      -- CP-element group 114: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/word_0/$exit
      -- CP-element group 114: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/word_0/ca
      -- 
    ca_3076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1148_store_0_ack_1, ack => convolution3D_CP_2151_elements(114)); -- 
    -- CP-element group 115:  branch  join  transition  place  output  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: 	76 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (10) 
      -- CP-element group 115: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161__exit__
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162__entry__
      -- CP-element group 115: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/$exit
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_dead_link/$entry
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_eval_test/$entry
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_eval_test/$exit
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_eval_test/branch_req
      -- CP-element group 115: 	 branch_block_stmt_720/R_exitcond23_1163_place
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_if_link/$entry
      -- CP-element group 115: 	 branch_block_stmt_720/if_stmt_1162_else_link/$entry
      -- 
    branch_req_3084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(115), ack => if_stmt_1162_branch_req_0); -- 
    convolution3D_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(114) & convolution3D_CP_2151_elements(76);
      gj_convolution3D_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  merge  transition  place  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	289 
    -- CP-element group 116:  members (13) 
      -- CP-element group 116: 	 branch_block_stmt_720/merge_stmt_1168__exit__
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xendx_xloopexit_forx_xend
      -- CP-element group 116: 	 branch_block_stmt_720/if_stmt_1162_if_link/$exit
      -- CP-element group 116: 	 branch_block_stmt_720/if_stmt_1162_if_link/if_choice_transition
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_720/merge_stmt_1168_PhiAck/dummy
      -- CP-element group 116: 	 branch_block_stmt_720/merge_stmt_1168_PhiAck/$exit
      -- CP-element group 116: 	 branch_block_stmt_720/merge_stmt_1168_PhiAck/$entry
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 116: 	 branch_block_stmt_720/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 116: 	 branch_block_stmt_720/merge_stmt_1168_PhiReqMerge
      -- 
    if_choice_transition_3089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1162_branch_ack_1, ack => convolution3D_CP_2151_elements(116)); -- 
    -- CP-element group 117:  fork  transition  place  input  output  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	284 
    -- CP-element group 117: 	285 
    -- CP-element group 117:  members (12) 
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/cr
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/rr
      -- CP-element group 117: 	 branch_block_stmt_720/if_stmt_1162_else_link/$exit
      -- CP-element group 117: 	 branch_block_stmt_720/if_stmt_1162_else_link/else_choice_transition
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/$entry
      -- CP-element group 117: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/$entry
      -- 
    else_choice_transition_3093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1162_branch_ack_0, ack => convolution3D_CP_2151_elements(117)); -- 
    cr_4342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(117), ack => type_cast_1005_inst_req_1); -- 
    rr_4337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(117), ack => type_cast_1005_inst_req_0); -- 
    -- CP-element group 118:  transition  input  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	289 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_sample_completed_
      -- CP-element group 118: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Sample/ra
      -- 
    ra_3107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => convolution3D_CP_2151_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	289 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	122 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_update_completed_
      -- CP-element group 119: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Update/ca
      -- 
    ca_3112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_1, ack => convolution3D_CP_2151_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	289 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Sample/$exit
      -- CP-element group 120: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Sample/ra
      -- 
    ra_3121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_0, ack => convolution3D_CP_2151_elements(120)); -- 
    -- CP-element group 121:  transition  input  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	289 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	122 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_update_completed_
      -- CP-element group 121: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Update/ca
      -- 
    ca_3126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1177_inst_ack_1, ack => convolution3D_CP_2151_elements(121)); -- 
    -- CP-element group 122:  branch  join  transition  place  output  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	119 
    -- CP-element group 122: 	121 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	123 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (10) 
      -- CP-element group 122: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199__exit__
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200__entry__
      -- CP-element group 122: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/$exit
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_dead_link/$entry
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_eval_test/$entry
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_eval_test/$exit
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_eval_test/branch_req
      -- CP-element group 122: 	 branch_block_stmt_720/R_cmp149340_1201_place
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_if_link/$entry
      -- CP-element group 122: 	 branch_block_stmt_720/if_stmt_1200_else_link/$entry
      -- 
    branch_req_3134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(122), ack => if_stmt_1200_branch_req_0); -- 
    convolution3D_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(119) & convolution3D_CP_2151_elements(121);
      gj_convolution3D_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	122 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	127 
    -- CP-element group 123: 	128 
    -- CP-element group 123: 	129 
    -- CP-element group 123: 	130 
    -- CP-element group 123: 	133 
    -- CP-element group 123: 	125 
    -- CP-element group 123: 	126 
    -- CP-element group 123:  members (33) 
      -- CP-element group 123: 	 branch_block_stmt_720/merge_stmt_1206__exit__
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280__entry__
      -- CP-element group 123: 	 branch_block_stmt_720/forx_xend_bbx_xnph_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/if_stmt_1200_if_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_720/if_stmt_1200_if_link/if_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_720/forx_xend_bbx_xnph
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_update_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_update_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_update_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_update_start_
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_720/merge_stmt_1206_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_720/merge_stmt_1206_PhiAck/dummy
      -- CP-element group 123: 	 branch_block_stmt_720/merge_stmt_1206_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_720/merge_stmt_1206_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_720/forx_xend_bbx_xnph_PhiReq/$exit
      -- 
    if_choice_transition_3139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1200_branch_ack_1, ack => convolution3D_CP_2151_elements(123)); -- 
    rr_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1221_inst_req_0); -- 
    cr_3161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1221_inst_req_1); -- 
    rr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3170_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1230_inst_req_0); -- 
    cr_3175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1230_inst_req_1); -- 
    rr_3184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1239_inst_req_0); -- 
    cr_3189_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3189_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1239_inst_req_1); -- 
    cr_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(123), ack => type_cast_1273_inst_req_1); -- 
    -- CP-element group 124:  transition  place  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	299 
    -- CP-element group 124:  members (6) 
      -- CP-element group 124: 	 branch_block_stmt_720/if_stmt_1200_else_link/$exit
      -- CP-element group 124: 	 branch_block_stmt_720/if_stmt_1200_else_link/else_choice_transition
      -- CP-element group 124: 	 branch_block_stmt_720/forx_xend_forx_xend203
      -- CP-element group 124: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$entry
      -- CP-element group 124: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/$entry
      -- CP-element group 124: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/$entry
      -- 
    else_choice_transition_3143_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1200_branch_ack_0, ack => convolution3D_CP_2151_elements(124)); -- 
    -- CP-element group 125:  transition  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Sample/ra
      -- 
    ra_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_0, ack => convolution3D_CP_2151_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	123 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	131 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1221_Update/ca
      -- 
    ca_3162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1221_inst_ack_1, ack => convolution3D_CP_2151_elements(126)); -- 
    -- CP-element group 127:  transition  input  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	123 
    -- CP-element group 127: successors 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Sample/ra
      -- 
    ra_3171_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_0, ack => convolution3D_CP_2151_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	123 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	131 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1230_Update/ca
      -- 
    ca_3176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1230_inst_ack_1, ack => convolution3D_CP_2151_elements(128)); -- 
    -- CP-element group 129:  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	123 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Sample/ra
      -- 
    ra_3185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_0, ack => convolution3D_CP_2151_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	123 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1239_Update/ca
      -- 
    ca_3190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1239_inst_ack_1, ack => convolution3D_CP_2151_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	128 
    -- CP-element group 131: 	130 
    -- CP-element group 131: 	126 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Sample/rr
      -- 
    rr_3198_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3198_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(131), ack => type_cast_1273_inst_req_0); -- 
    convolution3D_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(128) & convolution3D_CP_2151_elements(130) & convolution3D_CP_2151_elements(126);
      gj_convolution3D_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Sample/ra
      -- 
    ra_3199_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_0, ack => convolution3D_CP_2151_elements(132)); -- 
    -- CP-element group 133:  transition  place  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	123 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	290 
    -- CP-element group 133:  members (9) 
      -- CP-element group 133: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280__exit__
      -- CP-element group 133: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151
      -- CP-element group 133: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/$exit
      -- CP-element group 133: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_720/assign_stmt_1212_to_assign_stmt_1280/type_cast_1273_Update/ca
      -- CP-element group 133: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/$entry
      -- CP-element group 133: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/$entry
      -- CP-element group 133: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/$entry
      -- 
    ca_3204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1273_inst_ack_1, ack => convolution3D_CP_2151_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	295 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	173 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Sample/ack
      -- CP-element group 134: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_sample_complete
      -- 
    ack_3233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1295_index_offset_ack_0, ack => convolution3D_CP_2151_elements(134)); -- 
    -- CP-element group 135:  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	295 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (11) 
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_request/req
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_request/$entry
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_base_plus_offset/sum_rename_ack
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_base_plus_offset/sum_rename_req
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_base_plus_offset/$exit
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_base_plus_offset/$entry
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Update/ack
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_root_address_calculated
      -- CP-element group 135: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_offset_calculated
      -- 
    ack_3238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1295_index_offset_ack_1, ack => convolution3D_CP_2151_elements(135)); -- 
    req_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(135), ack => addr_of_1296_final_reg_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_request/ack
      -- CP-element group 136: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_request/$exit
      -- CP-element group 136: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_sample_completed_
      -- 
    ack_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1296_final_reg_ack_0, ack => convolution3D_CP_2151_elements(136)); -- 
    -- CP-element group 137:  fork  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	295 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	170 
    -- CP-element group 137:  members (19) 
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_plus_offset/$entry
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_addr_resize/base_resize_ack
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_word_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_addr_resize/base_resize_req
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_root_address_calculated
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_addr_resize/$entry
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_addr_resize/$exit
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_address_resized
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_plus_offset/$exit
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_complete/ack
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_complete/$exit
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_word_addrgen/root_register_ack
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_word_addrgen/root_register_req
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_word_addrgen/$exit
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_word_addrgen/$entry
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_plus_offset/sum_rename_ack
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_base_plus_offset/sum_rename_req
      -- CP-element group 137: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_update_completed_
      -- 
    ack_3253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1296_final_reg_ack_1, ack => convolution3D_CP_2151_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	295 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Update/cr
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_update_start_
      -- CP-element group 138: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_sample_completed_
      -- 
    ra_3262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1299_inst_ack_0, ack => convolution3D_CP_2151_elements(138)); -- 
    cr_3266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(138), ack => RPIPE_maxpool_input_pipe_1299_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_sample_start_
      -- 
    ca_3267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1299_inst_ack_1, ack => convolution3D_CP_2151_elements(139)); -- 
    rr_3275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(139), ack => type_cast_1303_inst_req_0); -- 
    rr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(139), ack => RPIPE_maxpool_input_pipe_1312_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Sample/ra
      -- CP-element group 140: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_sample_completed_
      -- 
    ra_3276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_0, ack => convolution3D_CP_2151_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	295 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	170 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Update/ca
      -- CP-element group 141: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Update/$exit
      -- 
    ca_3281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1303_inst_ack_1, ack => convolution3D_CP_2151_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Update/cr
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_update_start_
      -- CP-element group 142: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_sample_completed_
      -- 
    ra_3290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1312_inst_ack_0, ack => convolution3D_CP_2151_elements(142)); -- 
    cr_3294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(142), ack => RPIPE_maxpool_input_pipe_1312_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1312_update_completed_
      -- 
    ca_3295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1312_inst_ack_1, ack => convolution3D_CP_2151_elements(143)); -- 
    rr_3303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(143), ack => type_cast_1316_inst_req_0); -- 
    rr_3317_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3317_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(143), ack => RPIPE_maxpool_input_pipe_1330_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Sample/ra
      -- CP-element group 144: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_sample_completed_
      -- 
    ra_3304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_0, ack => convolution3D_CP_2151_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	295 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	170 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Update/ca
      -- CP-element group 145: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_update_completed_
      -- 
    ca_3309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1316_inst_ack_1, ack => convolution3D_CP_2151_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Update/cr
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_update_start_
      -- CP-element group 146: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_sample_completed_
      -- 
    ra_3318_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1330_inst_ack_0, ack => convolution3D_CP_2151_elements(146)); -- 
    cr_3322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(146), ack => RPIPE_maxpool_input_pipe_1330_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1330_update_completed_
      -- 
    ca_3323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1330_inst_ack_1, ack => convolution3D_CP_2151_elements(147)); -- 
    rr_3331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(147), ack => type_cast_1334_inst_req_0); -- 
    rr_3345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(147), ack => RPIPE_maxpool_input_pipe_1348_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Sample/ra
      -- CP-element group 148: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_sample_completed_
      -- 
    ra_3332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_0, ack => convolution3D_CP_2151_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	295 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	170 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Update/ca
      -- CP-element group 149: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_update_completed_
      -- 
    ca_3337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1334_inst_ack_1, ack => convolution3D_CP_2151_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Update/cr
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_update_start_
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Update/$entry
      -- 
    ra_3346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1348_inst_ack_0, ack => convolution3D_CP_2151_elements(150)); -- 
    cr_3350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(150), ack => RPIPE_maxpool_input_pipe_1348_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1348_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Sample/$entry
      -- 
    ca_3351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1348_inst_ack_1, ack => convolution3D_CP_2151_elements(151)); -- 
    rr_3359_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3359_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(151), ack => type_cast_1352_inst_req_0); -- 
    rr_3373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(151), ack => RPIPE_maxpool_input_pipe_1366_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Sample/ra
      -- CP-element group 152: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Sample/$exit
      -- 
    ra_3360_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1352_inst_ack_0, ack => convolution3D_CP_2151_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	295 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	170 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Update/ca
      -- CP-element group 153: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Update/$exit
      -- 
    ca_3365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1352_inst_ack_1, ack => convolution3D_CP_2151_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_update_start_
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Update/cr
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Sample/$exit
      -- 
    ra_3374_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1366_inst_ack_0, ack => convolution3D_CP_2151_elements(154)); -- 
    cr_3378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(154), ack => RPIPE_maxpool_input_pipe_1366_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1366_update_completed_
      -- 
    ca_3379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1366_inst_ack_1, ack => convolution3D_CP_2151_elements(155)); -- 
    rr_3387_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3387_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(155), ack => type_cast_1370_inst_req_0); -- 
    rr_3401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(155), ack => RPIPE_maxpool_input_pipe_1384_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Sample/ra
      -- CP-element group 156: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_sample_completed_
      -- 
    ra_3388_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_0, ack => convolution3D_CP_2151_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	295 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	170 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Update/ca
      -- CP-element group 157: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_update_completed_
      -- 
    ca_3393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1370_inst_ack_1, ack => convolution3D_CP_2151_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Update/cr
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_update_start_
      -- CP-element group 158: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_sample_completed_
      -- 
    ra_3402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_0, ack => convolution3D_CP_2151_elements(158)); -- 
    cr_3406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(158), ack => RPIPE_maxpool_input_pipe_1384_inst_req_1); -- 
    -- CP-element group 159:  fork  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159: 	162 
    -- CP-element group 159:  members (9) 
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Sample/rr
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1384_update_completed_
      -- 
    ca_3407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1384_inst_ack_1, ack => convolution3D_CP_2151_elements(159)); -- 
    rr_3415_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3415_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(159), ack => type_cast_1388_inst_req_0); -- 
    rr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(159), ack => RPIPE_maxpool_input_pipe_1402_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Sample/ra
      -- CP-element group 160: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_sample_completed_
      -- 
    ra_3416_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_0, ack => convolution3D_CP_2151_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	295 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	170 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Update/ca
      -- CP-element group 161: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_update_completed_
      -- 
    ca_3421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1388_inst_ack_1, ack => convolution3D_CP_2151_elements(161)); -- 
    -- CP-element group 162:  transition  input  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	159 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (6) 
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Sample/ra
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_sample_completed_
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Update/cr
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Sample/$exit
      -- CP-element group 162: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_update_start_
      -- 
    ra_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1402_inst_ack_0, ack => convolution3D_CP_2151_elements(162)); -- 
    cr_3434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(162), ack => RPIPE_maxpool_input_pipe_1402_inst_req_1); -- 
    -- CP-element group 163:  fork  transition  input  output  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	164 
    -- CP-element group 163: 	166 
    -- CP-element group 163:  members (9) 
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Update/$exit
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_Update/ca
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1402_update_completed_
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Sample/rr
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_sample_start_
      -- 
    ca_3435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1402_inst_ack_1, ack => convolution3D_CP_2151_elements(163)); -- 
    rr_3443_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3443_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(163), ack => type_cast_1406_inst_req_0); -- 
    rr_3457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(163), ack => RPIPE_maxpool_input_pipe_1420_inst_req_0); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	163 
    -- CP-element group 164: successors 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Sample/ra
      -- 
    ra_3444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_0, ack => convolution3D_CP_2151_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	295 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	170 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Update/ca
      -- CP-element group 165: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Update/$exit
      -- 
    ca_3449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1406_inst_ack_1, ack => convolution3D_CP_2151_elements(165)); -- 
    -- CP-element group 166:  transition  input  output  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	163 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	167 
    -- CP-element group 166:  members (6) 
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Update/cr
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Sample/ra
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Sample/$exit
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_update_start_
      -- CP-element group 166: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_sample_completed_
      -- 
    ra_3458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1420_inst_ack_0, ack => convolution3D_CP_2151_elements(166)); -- 
    cr_3462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(166), ack => RPIPE_maxpool_input_pipe_1420_inst_req_1); -- 
    -- CP-element group 167:  transition  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	166 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	168 
    -- CP-element group 167:  members (6) 
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Update/ca
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_Update/$exit
      -- CP-element group 167: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1420_update_completed_
      -- 
    ca_3463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1420_inst_ack_1, ack => convolution3D_CP_2151_elements(167)); -- 
    rr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3471_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(167), ack => type_cast_1424_inst_req_0); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	167 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Sample/ra
      -- CP-element group 168: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_sample_completed_
      -- 
    ra_3472_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1424_inst_ack_0, ack => convolution3D_CP_2151_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	295 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	170 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_update_completed_
      -- 
    ca_3477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1424_inst_ack_1, ack => convolution3D_CP_2151_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	137 
    -- CP-element group 170: 	141 
    -- CP-element group 170: 	145 
    -- CP-element group 170: 	149 
    -- CP-element group 170: 	153 
    -- CP-element group 170: 	157 
    -- CP-element group 170: 	161 
    -- CP-element group 170: 	165 
    -- CP-element group 170: 	169 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (9) 
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/word_0/rr
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/word_0/$entry
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/$entry
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/ptr_deref_1432_Split/split_ack
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/ptr_deref_1432_Split/split_req
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/ptr_deref_1432_Split/$exit
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/ptr_deref_1432_Split/$entry
      -- CP-element group 170: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/$entry
      -- 
    rr_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(170), ack => ptr_deref_1432_store_0_req_0); -- 
    convolution3D_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(137) & convolution3D_CP_2151_elements(141) & convolution3D_CP_2151_elements(145) & convolution3D_CP_2151_elements(149) & convolution3D_CP_2151_elements(153) & convolution3D_CP_2151_elements(157) & convolution3D_CP_2151_elements(161) & convolution3D_CP_2151_elements(165) & convolution3D_CP_2151_elements(169);
      gj_convolution3D_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	170 
    -- CP-element group 171: successors 
    -- CP-element group 171:  members (5) 
      -- CP-element group 171: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/word_0/ra
      -- CP-element group 171: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/word_0/$exit
      -- CP-element group 171: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/word_access_start/$exit
      -- CP-element group 171: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Sample/$exit
      -- 
    ra_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1432_store_0_ack_0, ack => convolution3D_CP_2151_elements(171)); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	295 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172:  members (5) 
      -- CP-element group 172: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/word_0/ca
      -- CP-element group 172: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/word_0/$exit
      -- CP-element group 172: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/$exit
      -- CP-element group 172: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/$exit
      -- 
    ca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1432_store_0_ack_1, ack => convolution3D_CP_2151_elements(172)); -- 
    -- CP-element group 173:  branch  join  transition  place  output  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: 	134 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	174 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (10) 
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_else_link/$entry
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_eval_test/branch_req
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_eval_test/$exit
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_eval_test/$entry
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_if_link/$entry
      -- CP-element group 173: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445__exit__
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446__entry__
      -- CP-element group 173: 	 branch_block_stmt_720/if_stmt_1446_dead_link/$entry
      -- CP-element group 173: 	 branch_block_stmt_720/R_exitcond22_1447_place
      -- CP-element group 173: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/$exit
      -- 
    branch_req_3535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(173), ack => if_stmt_1446_branch_req_0); -- 
    convolution3D_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(172) & convolution3D_CP_2151_elements(134);
      gj_convolution3D_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	173 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	177 
    -- CP-element group 174:  members (18) 
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Sample/rr
      -- CP-element group 174: 	 branch_block_stmt_720/if_stmt_1446_if_link/if_choice_transition
      -- CP-element group 174: 	 branch_block_stmt_720/if_stmt_1446_if_link/$exit
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/$entry
      -- CP-element group 174: 	 branch_block_stmt_720/merge_stmt_1452__exit__
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463__entry__
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_update_start_
      -- CP-element group 174: 	 branch_block_stmt_720/forx_xbody151_forx_xcond145x_xforx_xend203_crit_edge
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Update/cr
      -- CP-element group 174: 	 branch_block_stmt_720/merge_stmt_1452_PhiAck/dummy
      -- CP-element group 174: 	 branch_block_stmt_720/merge_stmt_1452_PhiAck/$exit
      -- CP-element group 174: 	 branch_block_stmt_720/merge_stmt_1452_PhiAck/$entry
      -- CP-element group 174: 	 branch_block_stmt_720/forx_xbody151_forx_xcond145x_xforx_xend203_crit_edge_PhiReq/$exit
      -- CP-element group 174: 	 branch_block_stmt_720/forx_xbody151_forx_xcond145x_xforx_xend203_crit_edge_PhiReq/$entry
      -- CP-element group 174: 	 branch_block_stmt_720/merge_stmt_1452_PhiReqMerge
      -- 
    if_choice_transition_3540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1446_branch_ack_1, ack => convolution3D_CP_2151_elements(174)); -- 
    rr_3557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(174), ack => type_cast_1462_inst_req_0); -- 
    cr_3562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(174), ack => type_cast_1462_inst_req_1); -- 
    -- CP-element group 175:  fork  transition  place  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	291 
    -- CP-element group 175: 	292 
    -- CP-element group 175:  members (12) 
      -- CP-element group 175: 	 branch_block_stmt_720/if_stmt_1446_else_link/$exit
      -- CP-element group 175: 	 branch_block_stmt_720/if_stmt_1446_else_link/else_choice_transition
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Update/cr
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/$entry
      -- CP-element group 175: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/$entry
      -- 
    else_choice_transition_3544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1446_branch_ack_0, ack => convolution3D_CP_2151_elements(175)); -- 
    cr_4419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(175), ack => type_cast_1289_inst_req_1); -- 
    rr_4414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(175), ack => type_cast_1289_inst_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Sample/ra
      -- CP-element group 176: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_sample_completed_
      -- 
    ra_3558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_0, ack => convolution3D_CP_2151_elements(176)); -- 
    -- CP-element group 177:  fork  transition  place  input  output  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	174 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	296 
    -- CP-element group 177: 	297 
    -- CP-element group 177:  members (15) 
      -- CP-element group 177: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463__exit__
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203
      -- CP-element group 177: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/$exit
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Update/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Sample/rr
      -- CP-element group 177: 	 branch_block_stmt_720/assign_stmt_1459_to_assign_stmt_1463/type_cast_1462_Update/ca
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/$entry
      -- CP-element group 177: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Update/cr
      -- 
    ca_3563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1462_inst_ack_1, ack => convolution3D_CP_2151_elements(177)); -- 
    rr_4457_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4457_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(177), ack => type_cast_1469_inst_req_0); -- 
    cr_4462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(177), ack => type_cast_1469_inst_req_1); -- 
    -- CP-element group 178:  transition  place  input  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	301 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	320 
    -- CP-element group 178:  members (5) 
      -- CP-element group 178: 	 branch_block_stmt_720/forx_xend203_ifx_xend
      -- CP-element group 178: 	 branch_block_stmt_720/if_stmt_1486_if_link/if_choice_transition
      -- CP-element group 178: 	 branch_block_stmt_720/if_stmt_1486_if_link/$exit
      -- CP-element group 178: 	 branch_block_stmt_720/forx_xend203_ifx_xend_PhiReq/$exit
      -- CP-element group 178: 	 branch_block_stmt_720/forx_xend203_ifx_xend_PhiReq/$entry
      -- 
    if_choice_transition_3579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1486_branch_ack_1, ack => convolution3D_CP_2151_elements(178)); -- 
    -- CP-element group 179:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	301 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	181 
    -- CP-element group 179: 	183 
    -- CP-element group 179:  members (21) 
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_720/forx_xend203_forx_xbodyx_xix_xpreheader
      -- CP-element group 179: 	 branch_block_stmt_720/merge_stmt_1492__exit__
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516__entry__
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Update/cr
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_update_start_
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_update_start_
      -- CP-element group 179: 	 branch_block_stmt_720/if_stmt_1486_else_link/else_choice_transition
      -- CP-element group 179: 	 branch_block_stmt_720/if_stmt_1486_else_link/$exit
      -- CP-element group 179: 	 branch_block_stmt_720/merge_stmt_1492_PhiAck/dummy
      -- CP-element group 179: 	 branch_block_stmt_720/merge_stmt_1492_PhiAck/$exit
      -- CP-element group 179: 	 branch_block_stmt_720/merge_stmt_1492_PhiAck/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/forx_xend203_forx_xbodyx_xix_xpreheader_PhiReq/$exit
      -- CP-element group 179: 	 branch_block_stmt_720/forx_xend203_forx_xbodyx_xix_xpreheader_PhiReq/$entry
      -- CP-element group 179: 	 branch_block_stmt_720/merge_stmt_1492_PhiReqMerge
      -- 
    else_choice_transition_3583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1486_branch_ack_0, ack => convolution3D_CP_2151_elements(179)); -- 
    cr_3601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(179), ack => type_cast_1511_inst_req_1); -- 
    rr_3596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(179), ack => type_cast_1511_inst_req_0); -- 
    cr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(179), ack => type_cast_1515_inst_req_1); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Sample/ra
      -- CP-element group 180: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_sample_completed_
      -- 
    ra_3597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_0, ack => convolution3D_CP_2151_elements(180)); -- 
    -- CP-element group 181:  transition  input  output  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	182 
    -- CP-element group 181:  members (6) 
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_Update/ca
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1511_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Sample/rr
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_sample_start_
      -- 
    ca_3602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_1, ack => convolution3D_CP_2151_elements(181)); -- 
    rr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(181), ack => type_cast_1515_inst_req_0); -- 
    -- CP-element group 182:  transition  input  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	181 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_sample_completed_
      -- 
    ra_3611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_0, ack => convolution3D_CP_2151_elements(182)); -- 
    -- CP-element group 183:  fork  transition  place  input  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	179 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	309 
    -- CP-element group 183: 	310 
    -- CP-element group 183:  members (11) 
      -- CP-element group 183: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516__exit__
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi
      -- CP-element group 183: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/$exit
      -- CP-element group 183: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_720/assign_stmt_1497_to_assign_stmt_1516/type_cast_1515_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$entry
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/$entry
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 183: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$entry
      -- 
    ca_3616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_1, ack => convolution3D_CP_2151_elements(183)); -- 
    -- CP-element group 184:  transition  input  output  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	315 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	185 
    -- CP-element group 184:  members (6) 
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_update_start_
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Update/cr
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Update/$entry
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Sample/ra
      -- CP-element group 184: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Sample/$exit
      -- 
    ra_3628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1535_inst_ack_0, ack => convolution3D_CP_2151_elements(184)); -- 
    cr_3632_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3632_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(184), ack => RPIPE_maxpool_input_pipe_1535_inst_req_1); -- 
    -- CP-element group 185:  transition  input  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	184 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	186 
    -- CP-element group 185:  members (6) 
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Update/ca
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_sample_start_
      -- 
    ca_3633_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_maxpool_input_pipe_1535_inst_ack_1, ack => convolution3D_CP_2151_elements(185)); -- 
    rr_3641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(185), ack => type_cast_1539_inst_req_0); -- 
    -- CP-element group 186:  transition  input  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	185 
    -- CP-element group 186: successors 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Sample/ra
      -- 
    ra_3642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_0, ack => convolution3D_CP_2151_elements(186)); -- 
    -- CP-element group 187:  branch  transition  place  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	315 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (13) 
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_eval_test/$exit
      -- CP-element group 187: 	 branch_block_stmt_720/R_exitcond2_1564_place
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_eval_test/branch_req
      -- CP-element group 187: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562__exit__
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563__entry__
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_dead_link/$entry
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_eval_test/$entry
      -- CP-element group 187: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/$exit
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_else_link/$entry
      -- CP-element group 187: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_720/if_stmt_1563_if_link/$entry
      -- 
    ca_3647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1539_inst_ack_1, ack => convolution3D_CP_2151_elements(187)); -- 
    branch_req_3655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(187), ack => if_stmt_1563_branch_req_0); -- 
    -- CP-element group 188:  fork  transition  place  input  output  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	316 
    -- CP-element group 188: 	317 
    -- CP-element group 188:  members (12) 
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit
      -- CP-element group 188: 	 branch_block_stmt_720/if_stmt_1563_if_link/if_choice_transition
      -- CP-element group 188: 	 branch_block_stmt_720/if_stmt_1563_if_link/$exit
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Update/cr
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Sample/rr
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Sample/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/$entry
      -- CP-element group 188: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$entry
      -- 
    if_choice_transition_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1563_branch_ack_1, ack => convolution3D_CP_2151_elements(188)); -- 
    cr_4594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(188), ack => type_cast_1573_inst_req_1); -- 
    rr_4589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(188), ack => type_cast_1573_inst_req_0); -- 
    -- CP-element group 189:  fork  transition  place  input  output  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	302 
    -- CP-element group 189: 	303 
    -- CP-element group 189: 	305 
    -- CP-element group 189: 	306 
    -- CP-element group 189:  members (20) 
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Update/cr
      -- CP-element group 189: 	 branch_block_stmt_720/if_stmt_1563_else_link/else_choice_transition
      -- CP-element group 189: 	 branch_block_stmt_720/if_stmt_1563_else_link/$exit
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/cr
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Sample/rr
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/$entry
      -- CP-element group 189: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/$entry
      -- 
    else_choice_transition_3664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1563_branch_ack_0, ack => convolution3D_CP_2151_elements(189)); -- 
    cr_4539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(189), ack => type_cast_1529_inst_req_1); -- 
    cr_4516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(189), ack => type_cast_1522_inst_req_1); -- 
    rr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(189), ack => type_cast_1522_inst_req_0); -- 
    rr_4534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(189), ack => type_cast_1529_inst_req_0); -- 
    -- CP-element group 190:  transition  input  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	319 
    -- CP-element group 190: successors 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Sample/ra
      -- 
    ra_3678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_0, ack => convolution3D_CP_2151_elements(190)); -- 
    -- CP-element group 191:  transition  input  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	319 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	196 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Update/ca
      -- 
    ca_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1577_inst_ack_1, ack => convolution3D_CP_2151_elements(191)); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	319 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	199 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_sample_complete
      -- CP-element group 192: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Sample/ack
      -- 
    ack_3709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1606_index_offset_ack_0, ack => convolution3D_CP_2151_elements(192)); -- 
    -- CP-element group 193:  transition  input  output  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	319 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (11) 
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_root_address_calculated
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_offset_calculated
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Update/ack
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_base_plus_offset/$entry
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_base_plus_offset/$exit
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_base_plus_offset/sum_rename_req
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_base_plus_offset/sum_rename_ack
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_request/$entry
      -- CP-element group 193: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_request/req
      -- 
    ack_3714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1606_index_offset_ack_1, ack => convolution3D_CP_2151_elements(193)); -- 
    req_3723_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3723_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(193), ack => addr_of_1607_final_reg_req_0); -- 
    -- CP-element group 194:  transition  input  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_request/$exit
      -- CP-element group 194: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_request/ack
      -- 
    ack_3724_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1607_final_reg_ack_0, ack => convolution3D_CP_2151_elements(194)); -- 
    -- CP-element group 195:  fork  transition  input  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	319 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (19) 
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_complete/$exit
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_complete/ack
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_word_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_root_address_calculated
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_address_resized
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_addr_resize/$entry
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_addr_resize/$exit
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_addr_resize/base_resize_req
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_addr_resize/base_resize_ack
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_plus_offset/$entry
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_plus_offset/$exit
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_plus_offset/sum_rename_req
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_base_plus_offset/sum_rename_ack
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_word_addrgen/$entry
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_word_addrgen/$exit
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_word_addrgen/root_register_req
      -- CP-element group 195: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_word_addrgen/root_register_ack
      -- 
    ack_3729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1607_final_reg_ack_1, ack => convolution3D_CP_2151_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	191 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196:  members (9) 
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/ptr_deref_1610_Split/$entry
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/ptr_deref_1610_Split/$exit
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/ptr_deref_1610_Split/split_req
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/ptr_deref_1610_Split/split_ack
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/$entry
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/word_0/$entry
      -- CP-element group 196: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/word_0/rr
      -- 
    rr_3767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(196), ack => ptr_deref_1610_store_0_req_0); -- 
    convolution3D_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(191) & convolution3D_CP_2151_elements(195);
      gj_convolution3D_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197:  members (5) 
      -- CP-element group 197: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_sample_completed_
      -- CP-element group 197: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/$exit
      -- CP-element group 197: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/$exit
      -- CP-element group 197: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/word_0/$exit
      -- CP-element group 197: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Sample/word_access_start/word_0/ra
      -- 
    ra_3768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1610_store_0_ack_0, ack => convolution3D_CP_2151_elements(197)); -- 
    -- CP-element group 198:  transition  input  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	319 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (5) 
      -- CP-element group 198: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_update_completed_
      -- CP-element group 198: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/$exit
      -- CP-element group 198: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/$exit
      -- CP-element group 198: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/word_0/$exit
      -- CP-element group 198: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/word_0/ca
      -- 
    ca_3779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1610_store_0_ack_1, ack => convolution3D_CP_2151_elements(198)); -- 
    -- CP-element group 199:  join  transition  place  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	192 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	320 
    -- CP-element group 199:  members (5) 
      -- CP-element group 199: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612__exit__
      -- CP-element group 199: 	 branch_block_stmt_720/getRemainingElementsx_xexit_ifx_xend
      -- CP-element group 199: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/$exit
      -- CP-element group 199: 	 branch_block_stmt_720/getRemainingElementsx_xexit_ifx_xend_PhiReq/$exit
      -- CP-element group 199: 	 branch_block_stmt_720/getRemainingElementsx_xexit_ifx_xend_PhiReq/$entry
      -- 
    convolution3D_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(192) & convolution3D_CP_2151_elements(198);
      gj_convolution3D_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	320 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Sample/cra
      -- 
    cra_3791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1617_call_ack_0, ack => convolution3D_CP_2151_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	320 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	208 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Update/cca
      -- 
    cca_3796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1617_call_ack_1, ack => convolution3D_CP_2151_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	320 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_update_start_
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Sample/ack
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Update/req
      -- 
    ack_3805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1618_inst_ack_0, ack => convolution3D_CP_2151_elements(202)); -- 
    req_3809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(202), ack => WPIPE_output_pipe_1618_inst_req_1); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Update/ack
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Sample/req
      -- 
    ack_3810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1618_inst_ack_1, ack => convolution3D_CP_2151_elements(203)); -- 
    req_3818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(203), ack => WPIPE_output_pipe_1621_inst_req_0); -- 
    -- CP-element group 204:  transition  input  output  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	205 
    -- CP-element group 204:  members (6) 
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_update_start_
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Sample/ack
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Update/req
      -- 
    ack_3819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1621_inst_ack_0, ack => convolution3D_CP_2151_elements(204)); -- 
    req_3823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(204), ack => WPIPE_output_pipe_1621_inst_req_1); -- 
    -- CP-element group 205:  transition  input  output  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	204 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (6) 
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1621_Update/ack
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_sample_start_
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Sample/$entry
      -- CP-element group 205: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Sample/req
      -- 
    ack_3824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1621_inst_ack_1, ack => convolution3D_CP_2151_elements(205)); -- 
    req_3832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(205), ack => WPIPE_output_pipe_1624_inst_req_0); -- 
    -- CP-element group 206:  transition  input  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (6) 
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_sample_completed_
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_update_start_
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Sample/$exit
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Sample/ack
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Update/$entry
      -- CP-element group 206: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Update/req
      -- 
    ack_3833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1624_inst_ack_0, ack => convolution3D_CP_2151_elements(206)); -- 
    req_3837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(206), ack => WPIPE_output_pipe_1624_inst_req_1); -- 
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_update_completed_
      -- CP-element group 207: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Update/$exit
      -- CP-element group 207: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1624_Update/ack
      -- 
    ack_3838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_1624_inst_ack_1, ack => convolution3D_CP_2151_elements(207)); -- 
    -- CP-element group 208:  join  fork  transition  place  output  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	201 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: 	210 
    -- CP-element group 208: 	211 
    -- CP-element group 208: 	212 
    -- CP-element group 208:  members (16) 
      -- CP-element group 208: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626__exit__
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669__entry__
      -- CP-element group 208: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/$exit
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/$entry
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_update_start_
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Update/cr
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_sample_start_
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_update_start_
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Sample/$entry
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Sample/rr
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Update/cr
      -- 
    rr_3849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(208), ack => type_cast_1642_inst_req_0); -- 
    cr_3854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(208), ack => type_cast_1642_inst_req_1); -- 
    rr_3863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(208), ack => type_cast_1663_inst_req_0); -- 
    cr_3868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(208), ack => type_cast_1663_inst_req_1); -- 
    convolution3D_cp_element_group_208: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_208"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(201) & convolution3D_CP_2151_elements(207);
      gj_convolution3D_cp_element_group_208 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(208), clk => clk, reset => reset); --
    end block;
    -- CP-element group 209:  transition  input  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_sample_completed_
      -- CP-element group 209: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Sample/$exit
      -- CP-element group 209: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Sample/ra
      -- 
    ra_3850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_0, ack => convolution3D_CP_2151_elements(209)); -- 
    -- CP-element group 210:  transition  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	208 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	213 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_update_completed_
      -- CP-element group 210: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Update/$exit
      -- CP-element group 210: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1642_Update/ca
      -- 
    ca_3855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1642_inst_ack_1, ack => convolution3D_CP_2151_elements(210)); -- 
    -- CP-element group 211:  transition  input  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	208 
    -- CP-element group 211: successors 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_sample_completed_
      -- CP-element group 211: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Sample/$exit
      -- CP-element group 211: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Sample/ra
      -- 
    ra_3864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_0, ack => convolution3D_CP_2151_elements(211)); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	208 
    -- CP-element group 212: successors 
    -- CP-element group 212: 	213 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_update_completed_
      -- CP-element group 212: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Update/$exit
      -- CP-element group 212: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/type_cast_1663_Update/ca
      -- 
    ca_3869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1663_inst_ack_1, ack => convolution3D_CP_2151_elements(212)); -- 
    -- CP-element group 213:  join  transition  place  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	210 
    -- CP-element group 213: 	212 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	321 
    -- CP-element group 213:  members (6) 
      -- CP-element group 213: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669__exit__
      -- CP-element group 213: 	 branch_block_stmt_720/ifx_xend_whilex_xbody
      -- CP-element group 213: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/$entry
      -- CP-element group 213: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/$entry
      -- CP-element group 213: 	 branch_block_stmt_720/assign_stmt_1633_to_assign_stmt_1669/$exit
      -- CP-element group 213: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/$entry
      -- 
    convolution3D_cp_element_group_213: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_213"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(210) & convolution3D_CP_2151_elements(212);
      gj_convolution3D_cp_element_group_213 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(213), clk => clk, reset => reset); --
    end block;
    -- CP-element group 214:  transition  input  output  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	326 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (6) 
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_update_start_
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Sample/$exit
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Sample/ack
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Update/$entry
      -- CP-element group 214: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Update/req
      -- 
    ack_3881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1685_inst_ack_0, ack => convolution3D_CP_2151_elements(214)); -- 
    req_3885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(214), ack => WPIPE_num_out_pipe_1685_inst_req_1); -- 
    -- CP-element group 215:  transition  input  output  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Update/$exit
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Update/ack
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_sample_start_
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Sample/$entry
      -- CP-element group 215: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Sample/req
      -- 
    ack_3886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1685_inst_ack_1, ack => convolution3D_CP_2151_elements(215)); -- 
    req_3894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(215), ack => WPIPE_num_out_pipe_1688_inst_req_0); -- 
    -- CP-element group 216:  transition  input  output  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	217 
    -- CP-element group 216:  members (6) 
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_update_start_
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Sample/ack
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Update/$entry
      -- CP-element group 216: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Update/req
      -- 
    ack_3895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1688_inst_ack_0, ack => convolution3D_CP_2151_elements(216)); -- 
    req_3899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(216), ack => WPIPE_num_out_pipe_1688_inst_req_1); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	216 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	222 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1688_Update/ack
      -- 
    ack_3900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_num_out_pipe_1688_inst_ack_1, ack => convolution3D_CP_2151_elements(217)); -- 
    -- CP-element group 218:  transition  input  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	326 
    -- CP-element group 218: successors 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_sample_completed_
      -- CP-element group 218: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Sample/$exit
      -- CP-element group 218: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Sample/cra
      -- 
    cra_3909_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 218_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1693_call_ack_0, ack => convolution3D_CP_2151_elements(218)); -- 
    -- CP-element group 219:  transition  input  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	326 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	222 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_update_completed_
      -- CP-element group 219: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Update/$exit
      -- CP-element group 219: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Update/cca
      -- 
    cca_3914_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1693_call_ack_1, ack => convolution3D_CP_2151_elements(219)); -- 
    -- CP-element group 220:  transition  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	326 
    -- CP-element group 220: successors 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Sample/cra
      -- 
    cra_3923_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1697_call_ack_0, ack => convolution3D_CP_2151_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	326 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	222 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Update/cca
      -- 
    cca_3928_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1697_call_ack_1, ack => convolution3D_CP_2151_elements(221)); -- 
    -- CP-element group 222:  branch  join  transition  place  output  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	221 
    -- CP-element group 222: 	217 
    -- CP-element group 222: 	219 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	223 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (10) 
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709__entry__
      -- CP-element group 222: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708__exit__
      -- CP-element group 222: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/$exit
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_dead_link/$entry
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_eval_test/$entry
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_eval_test/$exit
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_eval_test/branch_req
      -- CP-element group 222: 	 branch_block_stmt_720/R_exitcond_1710_place
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_if_link/$entry
      -- CP-element group 222: 	 branch_block_stmt_720/if_stmt_1709_else_link/$entry
      -- 
    branch_req_3936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(222), ack => if_stmt_1709_branch_req_0); -- 
    convolution3D_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(221) & convolution3D_CP_2151_elements(217) & convolution3D_CP_2151_elements(219);
      gj_convolution3D_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	222 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223: 	226 
    -- CP-element group 223: 	227 
    -- CP-element group 223:  members (21) 
      -- CP-element group 223: 	 branch_block_stmt_720/merge_stmt_1715__exit__
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724__entry__
      -- CP-element group 223: 	 branch_block_stmt_720/merge_stmt_1715_PhiReqMerge
      -- CP-element group 223: 	 branch_block_stmt_720/merge_stmt_1715_PhiAck/dummy
      -- CP-element group 223: 	 branch_block_stmt_720/merge_stmt_1715_PhiAck/$exit
      -- CP-element group 223: 	 branch_block_stmt_720/merge_stmt_1715_PhiAck/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/whilex_xbody_whilex_xend_PhiReq/$exit
      -- CP-element group 223: 	 branch_block_stmt_720/whilex_xbody_whilex_xend_PhiReq/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/if_stmt_1709_if_link/$exit
      -- CP-element group 223: 	 branch_block_stmt_720/if_stmt_1709_if_link/if_choice_transition
      -- CP-element group 223: 	 branch_block_stmt_720/whilex_xbody_whilex_xend
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_update_start_
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Sample/rr
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Update/cr
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_sample_start_
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Sample/$entry
      -- CP-element group 223: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Sample/rr
      -- 
    if_choice_transition_3941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1709_branch_ack_1, ack => convolution3D_CP_2151_elements(223)); -- 
    rr_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(223), ack => type_cast_1720_inst_req_0); -- 
    cr_3963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(223), ack => type_cast_1720_inst_req_1); -- 
    rr_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(223), ack => RPIPE_input_done_pipe_1723_inst_req_0); -- 
    -- CP-element group 224:  fork  transition  place  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	322 
    -- CP-element group 224: 	323 
    -- CP-element group 224:  members (12) 
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Update/cr
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Update/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Sample/rr
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Sample/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/if_stmt_1709_else_link/$exit
      -- CP-element group 224: 	 branch_block_stmt_720/if_stmt_1709_else_link/else_choice_transition
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/$entry
      -- CP-element group 224: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/$entry
      -- 
    else_choice_transition_3945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1709_branch_ack_0, ack => convolution3D_CP_2151_elements(224)); -- 
    cr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(224), ack => type_cast_1675_inst_req_1); -- 
    rr_4642_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4642_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(224), ack => type_cast_1675_inst_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Sample/$exit
      -- CP-element group 225: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Sample/ra
      -- 
    ra_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_0, ack => convolution3D_CP_2151_elements(225)); -- 
    -- CP-element group 226:  transition  input  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	223 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	229 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Update/$exit
      -- CP-element group 226: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/type_cast_1720_Update/ca
      -- 
    ca_3964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1720_inst_ack_1, ack => convolution3D_CP_2151_elements(226)); -- 
    -- CP-element group 227:  transition  input  output  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	223 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	228 
    -- CP-element group 227:  members (6) 
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_update_start_
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Sample/ra
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Update/cr
      -- 
    ra_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1723_inst_ack_0, ack => convolution3D_CP_2151_elements(227)); -- 
    cr_3977_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3977_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(227), ack => RPIPE_input_done_pipe_1723_inst_req_1); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	227 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/RPIPE_input_done_pipe_1723_Update/ca
      -- 
    ca_3978_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1723_inst_ack_1, ack => convolution3D_CP_2151_elements(228)); -- 
    -- CP-element group 229:  join  transition  place  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	226 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229:  members (7) 
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1728__entry__
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724__exit__
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1721_to_assign_stmt_1724/$exit
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1728/$entry
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Sample/rr
      -- 
    rr_3989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(229), ack => RPIPE_input_done_pipe_1727_inst_req_0); -- 
    convolution3D_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(226) & convolution3D_CP_2151_elements(228);
      gj_convolution3D_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  transition  input  output  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	231 
    -- CP-element group 230:  members (6) 
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_sample_completed_
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_update_start_
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Sample/$exit
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Sample/ra
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Update/cr
      -- 
    ra_3990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1727_inst_ack_0, ack => convolution3D_CP_2151_elements(230)); -- 
    cr_3994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(230), ack => RPIPE_input_done_pipe_1727_inst_req_1); -- 
    -- CP-element group 231:  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	230 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	232 
    -- CP-element group 231: 	233 
    -- CP-element group 231: 	235 
    -- CP-element group 231: 	236 
    -- CP-element group 231: 	237 
    -- CP-element group 231: 	238 
    -- CP-element group 231: 	239 
    -- CP-element group 231: 	242 
    -- CP-element group 231:  members (31) 
      -- CP-element group 231: 	 branch_block_stmt_720/assign_stmt_1728__exit__
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761__entry__
      -- CP-element group 231: 	 branch_block_stmt_720/assign_stmt_1728/$exit
      -- CP-element group 231: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_update_completed_
      -- CP-element group 231: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Update/$exit
      -- CP-element group 231: 	 branch_block_stmt_720/assign_stmt_1728/RPIPE_input_done_pipe_1727_Update/ca
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_update_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Sample/crr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Update/ccr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_update_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_update_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_sample_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_update_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Update/cr
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_update_start_
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Update/ccr
      -- 
    ca_3995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_1727_inst_ack_1, ack => convolution3D_CP_2151_elements(231)); -- 
    crr_4006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => call_stmt_1731_call_req_0); -- 
    ccr_4011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => call_stmt_1731_call_req_1); -- 
    cr_4025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => type_cast_1735_inst_req_1); -- 
    rr_4034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => type_cast_1744_inst_req_0); -- 
    cr_4039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => type_cast_1744_inst_req_1); -- 
    rr_4048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => type_cast_1748_inst_req_0); -- 
    cr_4053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => type_cast_1748_inst_req_1); -- 
    ccr_4067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(231), ack => call_stmt_1761_call_req_1); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	231 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Sample/cra
      -- 
    cra_4007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1731_call_ack_0, ack => convolution3D_CP_2151_elements(232)); -- 
    -- CP-element group 233:  transition  input  output  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	234 
    -- CP-element group 233:  members (6) 
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1731_Update/cca
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Sample/rr
      -- 
    cca_4012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1731_call_ack_1, ack => convolution3D_CP_2151_elements(233)); -- 
    rr_4020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(233), ack => type_cast_1735_inst_req_0); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	233 
    -- CP-element group 234: successors 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_sample_completed_
      -- CP-element group 234: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Sample/ra
      -- 
    ra_4021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1735_inst_ack_0, ack => convolution3D_CP_2151_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	231 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	243 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_update_completed_
      -- CP-element group 235: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1735_Update/ca
      -- 
    ca_4026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1735_inst_ack_1, ack => convolution3D_CP_2151_elements(235)); -- 
    -- CP-element group 236:  transition  input  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	231 
    -- CP-element group 236: successors 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Sample/ra
      -- 
    ra_4035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_0, ack => convolution3D_CP_2151_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	231 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	240 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1744_Update/ca
      -- 
    ca_4040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1744_inst_ack_1, ack => convolution3D_CP_2151_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	231 
    -- CP-element group 238: successors 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_sample_completed_
      -- CP-element group 238: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Sample/$exit
      -- CP-element group 238: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Sample/ra
      -- 
    ra_4049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_0, ack => convolution3D_CP_2151_elements(238)); -- 
    -- CP-element group 239:  transition  input  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	231 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_update_completed_
      -- CP-element group 239: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Update/$exit
      -- CP-element group 239: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/type_cast_1748_Update/ca
      -- 
    ca_4054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1748_inst_ack_1, ack => convolution3D_CP_2151_elements(239)); -- 
    -- CP-element group 240:  join  transition  output  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	237 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	241 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_sample_start_
      -- CP-element group 240: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Sample/$entry
      -- CP-element group 240: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Sample/crr
      -- 
    crr_4062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(240), ack => call_stmt_1761_call_req_0); -- 
    convolution3D_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(237) & convolution3D_CP_2151_elements(239);
      gj_convolution3D_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  transition  input  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	240 
    -- CP-element group 241: successors 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_sample_completed_
      -- CP-element group 241: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Sample/$exit
      -- CP-element group 241: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Sample/cra
      -- 
    cra_4063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1761_call_ack_0, ack => convolution3D_CP_2151_elements(241)); -- 
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	231 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	243 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_update_completed_
      -- CP-element group 242: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Update/$exit
      -- CP-element group 242: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/call_stmt_1761_Update/cca
      -- 
    cca_4068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1761_call_ack_1, ack => convolution3D_CP_2151_elements(242)); -- 
    -- CP-element group 243:  join  fork  transition  place  output  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	235 
    -- CP-element group 243: 	242 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243: 	245 
    -- CP-element group 243: 	246 
    -- CP-element group 243: 	247 
    -- CP-element group 243: 	248 
    -- CP-element group 243: 	249 
    -- CP-element group 243: 	250 
    -- CP-element group 243: 	251 
    -- CP-element group 243: 	252 
    -- CP-element group 243: 	253 
    -- CP-element group 243: 	254 
    -- CP-element group 243: 	255 
    -- CP-element group 243: 	256 
    -- CP-element group 243: 	257 
    -- CP-element group 243: 	258 
    -- CP-element group 243: 	259 
    -- CP-element group 243:  members (52) 
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860__entry__
      -- CP-element group 243: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761__exit__
      -- CP-element group 243: 	 branch_block_stmt_720/call_stmt_1731_to_call_stmt_1761/$exit
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Update/cr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_sample_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_update_start_
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Sample/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Sample/rr
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Update/cr
      -- 
    rr_4079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1765_inst_req_0); -- 
    cr_4084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1765_inst_req_1); -- 
    rr_4093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1775_inst_req_0); -- 
    cr_4098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1775_inst_req_1); -- 
    rr_4107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1785_inst_req_0); -- 
    cr_4112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1785_inst_req_1); -- 
    rr_4121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1795_inst_req_0); -- 
    cr_4126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1795_inst_req_1); -- 
    rr_4135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1805_inst_req_0); -- 
    cr_4140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1805_inst_req_1); -- 
    rr_4149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1815_inst_req_0); -- 
    cr_4154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1815_inst_req_1); -- 
    rr_4163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1825_inst_req_0); -- 
    cr_4168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1825_inst_req_1); -- 
    rr_4177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1835_inst_req_0); -- 
    cr_4182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(243), ack => type_cast_1835_inst_req_1); -- 
    convolution3D_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(235) & convolution3D_CP_2151_elements(242);
      gj_convolution3D_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  transition  input  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Sample/ra
      -- 
    ra_4080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1765_inst_ack_0, ack => convolution3D_CP_2151_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	280 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1765_Update/ca
      -- 
    ca_4085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1765_inst_ack_1, ack => convolution3D_CP_2151_elements(245)); -- 
    -- CP-element group 246:  transition  input  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	243 
    -- CP-element group 246: successors 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_sample_completed_
      -- CP-element group 246: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Sample/$exit
      -- CP-element group 246: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Sample/ra
      -- 
    ra_4094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 246_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1775_inst_ack_0, ack => convolution3D_CP_2151_elements(246)); -- 
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	243 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	277 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_update_completed_
      -- CP-element group 247: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Update/$exit
      -- CP-element group 247: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1775_Update/ca
      -- 
    ca_4099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1775_inst_ack_1, ack => convolution3D_CP_2151_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	243 
    -- CP-element group 248: successors 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Sample/ra
      -- 
    ra_4108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_0, ack => convolution3D_CP_2151_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	243 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	274 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1785_Update/ca
      -- 
    ca_4113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1785_inst_ack_1, ack => convolution3D_CP_2151_elements(249)); -- 
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	243 
    -- CP-element group 250: successors 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_sample_completed_
      -- CP-element group 250: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Sample/ra
      -- 
    ra_4122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_0, ack => convolution3D_CP_2151_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	243 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	271 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_update_completed_
      -- CP-element group 251: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1795_Update/ca
      -- 
    ca_4127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1795_inst_ack_1, ack => convolution3D_CP_2151_elements(251)); -- 
    -- CP-element group 252:  transition  input  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	243 
    -- CP-element group 252: successors 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Sample/ra
      -- 
    ra_4136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1805_inst_ack_0, ack => convolution3D_CP_2151_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	243 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	268 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1805_Update/ca
      -- 
    ca_4141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1805_inst_ack_1, ack => convolution3D_CP_2151_elements(253)); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	243 
    -- CP-element group 254: successors 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_sample_completed_
      -- CP-element group 254: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Sample/ra
      -- 
    ra_4150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_0, ack => convolution3D_CP_2151_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	243 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	265 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_update_completed_
      -- CP-element group 255: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1815_Update/ca
      -- 
    ca_4155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1815_inst_ack_1, ack => convolution3D_CP_2151_elements(255)); -- 
    -- CP-element group 256:  transition  input  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	243 
    -- CP-element group 256: successors 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Sample/ra
      -- 
    ra_4164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_0, ack => convolution3D_CP_2151_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	243 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	262 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1825_Update/ca
      -- 
    ca_4169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1825_inst_ack_1, ack => convolution3D_CP_2151_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	243 
    -- CP-element group 258: successors 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_sample_completed_
      -- CP-element group 258: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Sample/$exit
      -- CP-element group 258: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Sample/ra
      -- 
    ra_4178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_0, ack => convolution3D_CP_2151_elements(258)); -- 
    -- CP-element group 259:  transition  input  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	243 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_update_completed_
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Update/$exit
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/type_cast_1835_Update/ca
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_sample_start_
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Sample/$entry
      -- CP-element group 259: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Sample/req
      -- 
    ca_4183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1835_inst_ack_1, ack => convolution3D_CP_2151_elements(259)); -- 
    req_4191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(259), ack => WPIPE_maxpool_output_pipe_1837_inst_req_0); -- 
    -- CP-element group 260:  transition  input  output  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (6) 
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_update_start_
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Sample/ack
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Update/$entry
      -- CP-element group 260: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Update/req
      -- 
    ack_4192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1837_inst_ack_0, ack => convolution3D_CP_2151_elements(260)); -- 
    req_4196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(260), ack => WPIPE_maxpool_output_pipe_1837_inst_req_1); -- 
    -- CP-element group 261:  transition  input  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	262 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1837_Update/ack
      -- 
    ack_4197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1837_inst_ack_1, ack => convolution3D_CP_2151_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	257 
    -- CP-element group 262: 	261 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	263 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Sample/req
      -- 
    req_4205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(262), ack => WPIPE_maxpool_output_pipe_1840_inst_req_0); -- 
    convolution3D_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(257) & convolution3D_CP_2151_elements(261);
      gj_convolution3D_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  transition  input  output  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	262 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (6) 
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_update_start_
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Sample/ack
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Update/req
      -- 
    ack_4206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1840_inst_ack_0, ack => convolution3D_CP_2151_elements(263)); -- 
    req_4210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(263), ack => WPIPE_maxpool_output_pipe_1840_inst_req_1); -- 
    -- CP-element group 264:  transition  input  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	265 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1840_Update/ack
      -- 
    ack_4211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1840_inst_ack_1, ack => convolution3D_CP_2151_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	255 
    -- CP-element group 265: 	264 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_sample_start_
      -- CP-element group 265: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Sample/req
      -- 
    req_4219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(265), ack => WPIPE_maxpool_output_pipe_1843_inst_req_0); -- 
    convolution3D_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(255) & convolution3D_CP_2151_elements(264);
      gj_convolution3D_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  transition  input  output  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (6) 
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Update/req
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_sample_completed_
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_update_start_
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Sample/$exit
      -- CP-element group 266: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Sample/ack
      -- 
    ack_4220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 266_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1843_inst_ack_0, ack => convolution3D_CP_2151_elements(266)); -- 
    req_4224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(266), ack => WPIPE_maxpool_output_pipe_1843_inst_req_1); -- 
    -- CP-element group 267:  transition  input  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	268 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Update/ack
      -- CP-element group 267: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_Update/$exit
      -- CP-element group 267: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1843_update_completed_
      -- 
    ack_4225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1843_inst_ack_1, ack => convolution3D_CP_2151_elements(267)); -- 
    -- CP-element group 268:  join  transition  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	253 
    -- CP-element group 268: 	267 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	269 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Sample/req
      -- 
    req_4233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(268), ack => WPIPE_maxpool_output_pipe_1846_inst_req_0); -- 
    convolution3D_cp_element_group_268: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_268"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(253) & convolution3D_CP_2151_elements(267);
      gj_convolution3D_cp_element_group_268 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(268), clk => clk, reset => reset); --
    end block;
    -- CP-element group 269:  transition  input  output  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	268 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	270 
    -- CP-element group 269:  members (6) 
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_sample_completed_
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_update_start_
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Sample/$exit
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Update/req
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Update/$entry
      -- CP-element group 269: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Sample/ack
      -- 
    ack_4234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1846_inst_ack_0, ack => convolution3D_CP_2151_elements(269)); -- 
    req_4238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(269), ack => WPIPE_maxpool_output_pipe_1846_inst_req_1); -- 
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	269 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	271 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_update_completed_
      -- CP-element group 270: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Update/ack
      -- CP-element group 270: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1846_Update/$exit
      -- 
    ack_4239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1846_inst_ack_1, ack => convolution3D_CP_2151_elements(270)); -- 
    -- CP-element group 271:  join  transition  output  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	251 
    -- CP-element group 271: 	270 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Sample/$entry
      -- CP-element group 271: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_sample_start_
      -- CP-element group 271: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Sample/req
      -- 
    req_4247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(271), ack => WPIPE_maxpool_output_pipe_1849_inst_req_0); -- 
    convolution3D_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(251) & convolution3D_CP_2151_elements(270);
      gj_convolution3D_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  transition  input  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (6) 
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_update_start_
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Update/req
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Update/$entry
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Sample/ack
      -- CP-element group 272: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Sample/$exit
      -- 
    ack_4248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1849_inst_ack_0, ack => convolution3D_CP_2151_elements(272)); -- 
    req_4252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(272), ack => WPIPE_maxpool_output_pipe_1849_inst_req_1); -- 
    -- CP-element group 273:  transition  input  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	274 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Update/ack
      -- CP-element group 273: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1849_Update/$exit
      -- 
    ack_4253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1849_inst_ack_1, ack => convolution3D_CP_2151_elements(273)); -- 
    -- CP-element group 274:  join  transition  output  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	249 
    -- CP-element group 274: 	273 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	275 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Sample/req
      -- CP-element group 274: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_sample_start_
      -- 
    req_4261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(274), ack => WPIPE_maxpool_output_pipe_1852_inst_req_0); -- 
    convolution3D_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(249) & convolution3D_CP_2151_elements(273);
      gj_convolution3D_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  transition  input  output  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	274 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (6) 
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Sample/ack
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Update/req
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_update_start_
      -- CP-element group 275: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_sample_completed_
      -- 
    ack_4262_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1852_inst_ack_0, ack => convolution3D_CP_2151_elements(275)); -- 
    req_4266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(275), ack => WPIPE_maxpool_output_pipe_1852_inst_req_1); -- 
    -- CP-element group 276:  transition  input  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	277 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_update_completed_
      -- CP-element group 276: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1852_Update/ack
      -- 
    ack_4267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1852_inst_ack_1, ack => convolution3D_CP_2151_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	247 
    -- CP-element group 277: 	276 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	278 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Sample/req
      -- CP-element group 277: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Sample/$entry
      -- CP-element group 277: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_sample_start_
      -- 
    req_4275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(277), ack => WPIPE_maxpool_output_pipe_1855_inst_req_0); -- 
    convolution3D_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(247) & convolution3D_CP_2151_elements(276);
      gj_convolution3D_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  transition  input  output  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	277 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (6) 
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Sample/ack
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Sample/$exit
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_update_start_
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_sample_completed_
      -- CP-element group 278: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Update/req
      -- 
    ack_4276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1855_inst_ack_0, ack => convolution3D_CP_2151_elements(278)); -- 
    req_4280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(278), ack => WPIPE_maxpool_output_pipe_1855_inst_req_1); -- 
    -- CP-element group 279:  transition  input  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Update/$exit
      -- CP-element group 279: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_update_completed_
      -- CP-element group 279: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1855_Update/ack
      -- 
    ack_4281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1855_inst_ack_1, ack => convolution3D_CP_2151_elements(279)); -- 
    -- CP-element group 280:  join  transition  output  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	245 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Sample/req
      -- CP-element group 280: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Sample/$entry
      -- CP-element group 280: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_sample_start_
      -- 
    req_4289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(280), ack => WPIPE_maxpool_output_pipe_1858_inst_req_0); -- 
    convolution3D_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(245) & convolution3D_CP_2151_elements(279);
      gj_convolution3D_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  transition  input  output  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281:  members (6) 
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Update/req
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Update/$entry
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Sample/ack
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Sample/$exit
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_update_start_
      -- CP-element group 281: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_sample_completed_
      -- 
    ack_4290_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1858_inst_ack_0, ack => convolution3D_CP_2151_elements(281)); -- 
    req_4294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(281), ack => WPIPE_maxpool_output_pipe_1858_inst_req_1); -- 
    -- CP-element group 282:  transition  place  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282:  members (16) 
      -- CP-element group 282: 	 branch_block_stmt_720/merge_stmt_1862__exit__
      -- CP-element group 282: 	 branch_block_stmt_720/return__
      -- CP-element group 282: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860__exit__
      -- CP-element group 282: 	 branch_block_stmt_720/merge_stmt_1862_PhiReqMerge
      -- CP-element group 282: 	 $exit
      -- CP-element group 282: 	 branch_block_stmt_720/$exit
      -- CP-element group 282: 	 branch_block_stmt_720/branch_block_stmt_720__exit__
      -- CP-element group 282: 	 branch_block_stmt_720/merge_stmt_1862_PhiAck/$exit
      -- CP-element group 282: 	 branch_block_stmt_720/merge_stmt_1862_PhiAck/dummy
      -- CP-element group 282: 	 branch_block_stmt_720/return___PhiReq/$exit
      -- CP-element group 282: 	 branch_block_stmt_720/merge_stmt_1862_PhiAck/$entry
      -- CP-element group 282: 	 branch_block_stmt_720/return___PhiReq/$entry
      -- CP-element group 282: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Update/ack
      -- CP-element group 282: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_Update/$exit
      -- CP-element group 282: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/WPIPE_maxpool_output_pipe_1858_update_completed_
      -- CP-element group 282: 	 branch_block_stmt_720/assign_stmt_1766_to_assign_stmt_1860/$exit
      -- 
    ack_4295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_1858_inst_ack_1, ack => convolution3D_CP_2151_elements(282)); -- 
    -- CP-element group 283:  transition  output  delay-element  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	75 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	287 
    -- CP-element group 283:  members (5) 
      -- CP-element group 283: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_req
      -- CP-element group 283: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1003_konst_delay_trans
      -- CP-element group 283: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/$exit
      -- CP-element group 283: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/phi_stmt_999/$exit
      -- CP-element group 283: 	 branch_block_stmt_720/bbx_xnph345_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_999_req_4318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_999_req_4318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(283), ack => phi_stmt_999_req_0); -- 
    -- Element group convolution3D_CP_2151_elements(283) is a control-delay.
    cp_element_283_delay: control_delay_element  generic map(name => " 283_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(75), ack => convolution3D_CP_2151_elements(283), clk => clk, reset =>reset);
    -- CP-element group 284:  transition  input  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	117 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	286 
    -- CP-element group 284:  members (2) 
      -- CP-element group 284: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/ra
      -- CP-element group 284: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Sample/$exit
      -- 
    ra_4338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_0, ack => convolution3D_CP_2151_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	117 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	286 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/Update/ca
      -- 
    ca_4343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1005_inst_ack_1, ack => convolution3D_CP_2151_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	284 
    -- CP-element group 286: 	285 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (6) 
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_req
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/SplitProtocol/$exit
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/type_cast_1005/$exit
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/phi_stmt_999_sources/$exit
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/phi_stmt_999/$exit
      -- CP-element group 286: 	 branch_block_stmt_720/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    phi_stmt_999_req_4344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_999_req_4344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(286), ack => phi_stmt_999_req_1); -- 
    convolution3D_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(284) & convolution3D_CP_2151_elements(285);
      gj_convolution3D_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  merge  transition  place  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	283 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (2) 
      -- CP-element group 287: 	 branch_block_stmt_720/merge_stmt_998_PhiAck/$entry
      -- CP-element group 287: 	 branch_block_stmt_720/merge_stmt_998_PhiReqMerge
      -- 
    convolution3D_CP_2151_elements(287) <= OrReduce(convolution3D_CP_2151_elements(283) & convolution3D_CP_2151_elements(286));
    -- CP-element group 288:  fork  transition  place  input  output  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	83 
    -- CP-element group 288: 	87 
    -- CP-element group 288: 	91 
    -- CP-element group 288: 	95 
    -- CP-element group 288: 	99 
    -- CP-element group 288: 	103 
    -- CP-element group 288: 	107 
    -- CP-element group 288: 	111 
    -- CP-element group 288: 	114 
    -- CP-element group 288: 	76 
    -- CP-element group 288: 	77 
    -- CP-element group 288: 	79 
    -- CP-element group 288: 	80 
    -- CP-element group 288:  members (56) 
      -- CP-element group 288: 	 branch_block_stmt_720/merge_stmt_998__exit__
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161__entry__
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_resized_1
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_scaled_1
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_computed_1
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_resize_1/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_resize_1/$exit
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_resize_1/index_resize_req
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_resize_1/index_resize_ack
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_scale_1/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_scale_1/$exit
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_scale_1/scale_rename_req
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_index_scale_1/scale_rename_ack
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_update_start
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Sample/req
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/array_obj_ref_1011_final_index_sum_regn_Update/req
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_complete/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/addr_of_1012_complete/req
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_sample_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Sample/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/RPIPE_maxpool_input_pipe_1015_Sample/rr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1019_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1032_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1050_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1068_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1086_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1104_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1122_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/type_cast_1140_Update/cr
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_update_start_
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/word_0/$entry
      -- CP-element group 288: 	 branch_block_stmt_720/assign_stmt_1013_to_assign_stmt_1161/ptr_deref_1148_Update/word_access_complete/word_0/cr
      -- CP-element group 288: 	 branch_block_stmt_720/merge_stmt_998_PhiAck/$exit
      -- CP-element group 288: 	 branch_block_stmt_720/merge_stmt_998_PhiAck/phi_stmt_999_ack
      -- 
    phi_stmt_999_ack_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_999_ack_0, ack => convolution3D_CP_2151_elements(288)); -- 
    req_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => array_obj_ref_1011_index_offset_req_0); -- 
    req_2786_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2786_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => array_obj_ref_1011_index_offset_req_1); -- 
    req_2801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => addr_of_1012_final_reg_req_1); -- 
    rr_2810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => RPIPE_maxpool_input_pipe_1015_inst_req_0); -- 
    cr_2829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1019_inst_req_1); -- 
    cr_2857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1032_inst_req_1); -- 
    cr_2885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1050_inst_req_1); -- 
    cr_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1068_inst_req_1); -- 
    cr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1086_inst_req_1); -- 
    cr_2969_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2969_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1104_inst_req_1); -- 
    cr_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1122_inst_req_1); -- 
    cr_3025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => type_cast_1140_inst_req_1); -- 
    cr_3075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(288), ack => ptr_deref_1148_store_0_req_1); -- 
    -- CP-element group 289:  merge  fork  transition  place  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	116 
    -- CP-element group 289: 	73 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	118 
    -- CP-element group 289: 	119 
    -- CP-element group 289: 	120 
    -- CP-element group 289: 	121 
    -- CP-element group 289:  members (19) 
      -- CP-element group 289: 	 branch_block_stmt_720/merge_stmt_1170__exit__
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199__entry__
      -- CP-element group 289: 	 branch_block_stmt_720/merge_stmt_1170_PhiAck/dummy
      -- CP-element group 289: 	 branch_block_stmt_720/merge_stmt_1170_PhiAck/$exit
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_update_start_
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1173_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_sample_start_
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_update_start_
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Update/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/assign_stmt_1174_to_assign_stmt_1199/type_cast_1177_Update/cr
      -- CP-element group 289: 	 branch_block_stmt_720/merge_stmt_1170_PhiAck/$entry
      -- CP-element group 289: 	 branch_block_stmt_720/merge_stmt_1170_PhiReqMerge
      -- 
    rr_3106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(289), ack => type_cast_1173_inst_req_0); -- 
    cr_3111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(289), ack => type_cast_1173_inst_req_1); -- 
    rr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(289), ack => type_cast_1177_inst_req_0); -- 
    cr_3125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(289), ack => type_cast_1177_inst_req_1); -- 
    convolution3D_CP_2151_elements(289) <= OrReduce(convolution3D_CP_2151_elements(116) & convolution3D_CP_2151_elements(73));
    -- CP-element group 290:  transition  output  delay-element  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	133 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	294 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_req
      -- CP-element group 290: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1287_konst_delay_trans
      -- CP-element group 290: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/phi_stmt_1283/$exit
      -- CP-element group 290: 	 branch_block_stmt_720/bbx_xnph_forx_xbody151_PhiReq/$exit
      -- 
    phi_stmt_1283_req_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1283_req_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(290), ack => phi_stmt_1283_req_0); -- 
    -- Element group convolution3D_CP_2151_elements(290) is a control-delay.
    cp_element_290_delay: control_delay_element  generic map(name => " 290_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(133), ack => convolution3D_CP_2151_elements(290), clk => clk, reset =>reset);
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	175 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (2) 
      -- CP-element group 291: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Sample/ra
      -- CP-element group 291: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Sample/$exit
      -- 
    ra_4415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_0, ack => convolution3D_CP_2151_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	175 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Update/ca
      -- CP-element group 292: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/Update/$exit
      -- 
    ca_4420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1289_inst_ack_1, ack => convolution3D_CP_2151_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_req
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/SplitProtocol/$exit
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/type_cast_1289/$exit
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/phi_stmt_1283_sources/$exit
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/phi_stmt_1283/$exit
      -- CP-element group 293: 	 branch_block_stmt_720/forx_xbody151_forx_xbody151_PhiReq/$exit
      -- 
    phi_stmt_1283_req_4421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1283_req_4421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(293), ack => phi_stmt_1283_req_1); -- 
    convolution3D_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(291) & convolution3D_CP_2151_elements(292);
      gj_convolution3D_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  merge  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	290 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_720/merge_stmt_1282_PhiAck/$entry
      -- CP-element group 294: 	 branch_block_stmt_720/merge_stmt_1282_PhiReqMerge
      -- 
    convolution3D_CP_2151_elements(294) <= OrReduce(convolution3D_CP_2151_elements(290) & convolution3D_CP_2151_elements(293));
    -- CP-element group 295:  fork  transition  place  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	137 
    -- CP-element group 295: 	138 
    -- CP-element group 295: 	141 
    -- CP-element group 295: 	145 
    -- CP-element group 295: 	149 
    -- CP-element group 295: 	153 
    -- CP-element group 295: 	157 
    -- CP-element group 295: 	161 
    -- CP-element group 295: 	165 
    -- CP-element group 295: 	169 
    -- CP-element group 295: 	172 
    -- CP-element group 295: 	134 
    -- CP-element group 295: 	135 
    -- CP-element group 295:  members (56) 
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_scale_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/merge_stmt_1282__exit__
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445__entry__
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1352_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_update_start
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_scale_1/scale_rename_ack
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1334_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/word_0/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/RPIPE_maxpool_input_pipe_1299_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1388_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_complete/req
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1424_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/ptr_deref_1432_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_scale_1/scale_rename_req
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_resize_1/index_resize_ack
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_scale_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1370_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1406_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1316_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_resize_1/index_resize_req
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_resize_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_final_index_sum_regn_Update/req
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_resize_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/type_cast_1303_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/$entry
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/addr_of_1296_update_start_
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_resized_1
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_scaled_1
      -- CP-element group 295: 	 branch_block_stmt_720/assign_stmt_1297_to_assign_stmt_1445/array_obj_ref_1295_index_computed_1
      -- CP-element group 295: 	 branch_block_stmt_720/merge_stmt_1282_PhiAck/phi_stmt_1283_ack
      -- CP-element group 295: 	 branch_block_stmt_720/merge_stmt_1282_PhiAck/$exit
      -- 
    phi_stmt_1283_ack_4426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1283_ack_0, ack => convolution3D_CP_2151_elements(295)); -- 
    cr_3420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1388_inst_req_1); -- 
    cr_3336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1334_inst_req_1); -- 
    rr_3261_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3261_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => RPIPE_maxpool_input_pipe_1299_inst_req_0); -- 
    req_3232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => array_obj_ref_1295_index_offset_req_0); -- 
    cr_3364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1352_inst_req_1); -- 
    cr_3476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1424_inst_req_1); -- 
    cr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => ptr_deref_1432_store_0_req_1); -- 
    req_3252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => addr_of_1296_final_reg_req_1); -- 
    cr_3392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1370_inst_req_1); -- 
    cr_3308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1316_inst_req_1); -- 
    cr_3448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1406_inst_req_1); -- 
    req_3237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => array_obj_ref_1295_index_offset_req_1); -- 
    cr_3280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(295), ack => type_cast_1303_inst_req_1); -- 
    -- CP-element group 296:  transition  input  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	177 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	298 
    -- CP-element group 296:  members (2) 
      -- CP-element group 296: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Sample/ra
      -- CP-element group 296: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Sample/$exit
      -- 
    ra_4458_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_0, ack => convolution3D_CP_2151_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	177 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	298 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/Update/ca
      -- 
    ca_4463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1469_inst_ack_1, ack => convolution3D_CP_2151_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	296 
    -- CP-element group 298: 	297 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (6) 
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/SplitProtocol/$exit
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1469/$exit
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$exit
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/$exit
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/$exit
      -- CP-element group 298: 	 branch_block_stmt_720/forx_xcond145x_xforx_xend203_crit_edge_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_req
      -- 
    phi_stmt_1466_req_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1466_req_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(298), ack => phi_stmt_1466_req_0); -- 
    convolution3D_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(296) & convolution3D_CP_2151_elements(297);
      gj_convolution3D_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  transition  output  delay-element  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	124 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (5) 
      -- CP-element group 299: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_req
      -- CP-element group 299: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/type_cast_1472_konst_delay_trans
      -- CP-element group 299: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/phi_stmt_1466_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/phi_stmt_1466/$exit
      -- CP-element group 299: 	 branch_block_stmt_720/forx_xend_forx_xend203_PhiReq/$exit
      -- 
    phi_stmt_1466_req_4475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1466_req_4475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(299), ack => phi_stmt_1466_req_1); -- 
    -- Element group convolution3D_CP_2151_elements(299) is a control-delay.
    cp_element_299_delay: control_delay_element  generic map(name => " 299_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(124), ack => convolution3D_CP_2151_elements(299), clk => clk, reset =>reset);
    -- CP-element group 300:  merge  transition  place  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_720/merge_stmt_1465_PhiReqMerge
      -- CP-element group 300: 	 branch_block_stmt_720/merge_stmt_1465_PhiAck/$entry
      -- 
    convolution3D_CP_2151_elements(300) <= OrReduce(convolution3D_CP_2151_elements(298) & convolution3D_CP_2151_elements(299));
    -- CP-element group 301:  branch  transition  place  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	178 
    -- CP-element group 301: 	179 
    -- CP-element group 301:  members (15) 
      -- CP-element group 301: 	 branch_block_stmt_720/R_tobool_1487_place
      -- CP-element group 301: 	 branch_block_stmt_720/merge_stmt_1465__exit__
      -- CP-element group 301: 	 branch_block_stmt_720/assign_stmt_1479_to_assign_stmt_1485__entry__
      -- CP-element group 301: 	 branch_block_stmt_720/assign_stmt_1479_to_assign_stmt_1485__exit__
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486__entry__
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_dead_link/$entry
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_else_link/$entry
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_if_link/$entry
      -- CP-element group 301: 	 branch_block_stmt_720/assign_stmt_1479_to_assign_stmt_1485/$exit
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_eval_test/branch_req
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_eval_test/$exit
      -- CP-element group 301: 	 branch_block_stmt_720/if_stmt_1486_eval_test/$entry
      -- CP-element group 301: 	 branch_block_stmt_720/assign_stmt_1479_to_assign_stmt_1485/$entry
      -- CP-element group 301: 	 branch_block_stmt_720/merge_stmt_1465_PhiAck/phi_stmt_1466_ack
      -- CP-element group 301: 	 branch_block_stmt_720/merge_stmt_1465_PhiAck/$exit
      -- 
    phi_stmt_1466_ack_4480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1466_ack_0, ack => convolution3D_CP_2151_elements(301)); -- 
    branch_req_3574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(301), ack => if_stmt_1486_branch_req_0); -- 
    -- CP-element group 302:  transition  input  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	189 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (2) 
      -- CP-element group 302: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/ra
      -- CP-element group 302: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Sample/$exit
      -- 
    ra_4512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 302_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_0, ack => convolution3D_CP_2151_elements(302)); -- 
    -- CP-element group 303:  transition  input  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	189 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	304 
    -- CP-element group 303:  members (2) 
      -- CP-element group 303: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/ca
      -- CP-element group 303: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/Update/$exit
      -- 
    ca_4517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1522_inst_ack_1, ack => convolution3D_CP_2151_elements(303)); -- 
    -- CP-element group 304:  join  transition  output  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: 	303 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	308 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_req
      -- CP-element group 304: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/SplitProtocol/$exit
      -- CP-element group 304: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1522/$exit
      -- CP-element group 304: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$exit
      -- CP-element group 304: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1519/$exit
      -- 
    phi_stmt_1519_req_4518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1519_req_4518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(304), ack => phi_stmt_1519_req_0); -- 
    convolution3D_cp_element_group_304: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_304"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(302) & convolution3D_CP_2151_elements(303);
      gj_convolution3D_cp_element_group_304 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(304), clk => clk, reset => reset); --
    end block;
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	189 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Sample/ra
      -- CP-element group 305: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Sample/$exit
      -- 
    ra_4535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_0, ack => convolution3D_CP_2151_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	189 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Update/ca
      -- CP-element group 306: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/Update/$exit
      -- 
    ca_4540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1529_inst_ack_1, ack => convolution3D_CP_2151_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (5) 
      -- CP-element group 307: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- CP-element group 307: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/$exit
      -- CP-element group 307: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1529/$exit
      -- 
    phi_stmt_1526_req_4541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_4541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(307), ack => phi_stmt_1526_req_0); -- 
    convolution3D_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(305) & convolution3D_CP_2151_elements(306);
      gj_convolution3D_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  join  transition  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	304 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	312 
    -- CP-element group 308:  members (1) 
      -- CP-element group 308: 	 branch_block_stmt_720/forx_xbodyx_xi_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_308: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_308"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(304) & convolution3D_CP_2151_elements(307);
      gj_convolution3D_cp_element_group_308 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(308), clk => clk, reset => reset); --
    end block;
    -- CP-element group 309:  transition  output  delay-element  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	183 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (4) 
      -- CP-element group 309: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/$exit
      -- CP-element group 309: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/$exit
      -- CP-element group 309: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_req
      -- CP-element group 309: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1519/phi_stmt_1519_sources/type_cast_1525_konst_delay_trans
      -- 
    phi_stmt_1519_req_4552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1519_req_4552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(309), ack => phi_stmt_1519_req_1); -- 
    -- Element group convolution3D_CP_2151_elements(309) is a control-delay.
    cp_element_309_delay: control_delay_element  generic map(name => " 309_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(183), ack => convolution3D_CP_2151_elements(309), clk => clk, reset =>reset);
    -- CP-element group 310:  transition  output  delay-element  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	183 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	311 
    -- CP-element group 310:  members (4) 
      -- CP-element group 310: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_req
      -- CP-element group 310: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/type_cast_1532_konst_delay_trans
      -- CP-element group 310: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/phi_stmt_1526_sources/$exit
      -- CP-element group 310: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/phi_stmt_1526/$exit
      -- 
    phi_stmt_1526_req_4560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1526_req_4560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(310), ack => phi_stmt_1526_req_1); -- 
    -- Element group convolution3D_CP_2151_elements(310) is a control-delay.
    cp_element_310_delay: control_delay_element  generic map(name => " 310_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(183), ack => convolution3D_CP_2151_elements(310), clk => clk, reset =>reset);
    -- CP-element group 311:  join  transition  bypass 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	310 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	312 
    -- CP-element group 311:  members (1) 
      -- CP-element group 311: 	 branch_block_stmt_720/forx_xbodyx_xix_xpreheader_forx_xbodyx_xi_PhiReq/$exit
      -- 
    convolution3D_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(309) & convolution3D_CP_2151_elements(310);
      gj_convolution3D_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  merge  fork  transition  place  bypass 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	308 
    -- CP-element group 312: 	311 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	313 
    -- CP-element group 312: 	314 
    -- CP-element group 312:  members (2) 
      -- CP-element group 312: 	 branch_block_stmt_720/merge_stmt_1518_PhiReqMerge
      -- CP-element group 312: 	 branch_block_stmt_720/merge_stmt_1518_PhiAck/$entry
      -- 
    convolution3D_CP_2151_elements(312) <= OrReduce(convolution3D_CP_2151_elements(308) & convolution3D_CP_2151_elements(311));
    -- CP-element group 313:  transition  input  bypass 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	312 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (1) 
      -- CP-element group 313: 	 branch_block_stmt_720/merge_stmt_1518_PhiAck/phi_stmt_1519_ack
      -- 
    phi_stmt_1519_ack_4565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1519_ack_0, ack => convolution3D_CP_2151_elements(313)); -- 
    -- CP-element group 314:  transition  input  bypass 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	312 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	315 
    -- CP-element group 314:  members (1) 
      -- CP-element group 314: 	 branch_block_stmt_720/merge_stmt_1518_PhiAck/phi_stmt_1526_ack
      -- 
    phi_stmt_1526_ack_4566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 314_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1526_ack_0, ack => convolution3D_CP_2151_elements(314)); -- 
    -- CP-element group 315:  join  fork  transition  place  output  bypass 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	314 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	184 
    -- CP-element group 315: 	187 
    -- CP-element group 315:  members (10) 
      -- CP-element group 315: 	 branch_block_stmt_720/merge_stmt_1518__exit__
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562__entry__
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_sample_start_
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Sample/rr
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/$entry
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/RPIPE_maxpool_input_pipe_1535_Sample/$entry
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_update_start_
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Update/cr
      -- CP-element group 315: 	 branch_block_stmt_720/assign_stmt_1536_to_assign_stmt_1562/type_cast_1539_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_720/merge_stmt_1518_PhiAck/$exit
      -- 
    rr_3627_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3627_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(315), ack => RPIPE_maxpool_input_pipe_1535_inst_req_0); -- 
    cr_3646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(315), ack => type_cast_1539_inst_req_1); -- 
    convolution3D_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(313) & convolution3D_CP_2151_elements(314);
      gj_convolution3D_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  transition  input  bypass 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	188 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	318 
    -- CP-element group 316:  members (2) 
      -- CP-element group 316: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Sample/$exit
      -- 
    ra_4590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1573_inst_ack_0, ack => convolution3D_CP_2151_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	188 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	318 
    -- CP-element group 317:  members (2) 
      -- CP-element group 317: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Update/ca
      -- CP-element group 317: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/Update/$exit
      -- 
    ca_4595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1573_inst_ack_1, ack => convolution3D_CP_2151_elements(317)); -- 
    -- CP-element group 318:  join  transition  place  output  bypass 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	316 
    -- CP-element group 318: 	317 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	319 
    -- CP-element group 318:  members (8) 
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_req
      -- CP-element group 318: 	 branch_block_stmt_720/merge_stmt_1569_PhiReqMerge
      -- CP-element group 318: 	 branch_block_stmt_720/merge_stmt_1569_PhiAck/$entry
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/SplitProtocol/$exit
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/type_cast_1573/$exit
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/phi_stmt_1570_sources/$exit
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/phi_stmt_1570/$exit
      -- CP-element group 318: 	 branch_block_stmt_720/forx_xbodyx_xi_getRemainingElementsx_xexit_PhiReq/$exit
      -- 
    phi_stmt_1570_req_4596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1570_req_4596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(318), ack => phi_stmt_1570_req_0); -- 
    convolution3D_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(316) & convolution3D_CP_2151_elements(317);
      gj_convolution3D_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	318 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	190 
    -- CP-element group 319: 	191 
    -- CP-element group 319: 	192 
    -- CP-element group 319: 	193 
    -- CP-element group 319: 	195 
    -- CP-element group 319: 	198 
    -- CP-element group 319:  members (35) 
      -- CP-element group 319: 	 branch_block_stmt_720/merge_stmt_1569__exit__
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612__entry__
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_sample_start_
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_update_start_
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Sample/rr
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/type_cast_1577_Update/cr
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_update_start_
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_resized_1
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_scaled_1
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_computed_1
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_resize_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_resize_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_resize_1/index_resize_req
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_resize_1/index_resize_ack
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_scale_1/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_scale_1/$exit
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_scale_1/scale_rename_req
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_index_scale_1/scale_rename_ack
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_update_start
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Sample/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Sample/req
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/array_obj_ref_1606_final_index_sum_regn_Update/req
      -- CP-element group 319: 	 branch_block_stmt_720/merge_stmt_1569_PhiAck/phi_stmt_1570_ack
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/merge_stmt_1569_PhiAck/$exit
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/addr_of_1607_complete/req
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_update_start_
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/word_0/$entry
      -- CP-element group 319: 	 branch_block_stmt_720/assign_stmt_1578_to_assign_stmt_1612/ptr_deref_1610_Update/word_access_complete/word_0/cr
      -- 
    phi_stmt_1570_ack_4601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1570_ack_0, ack => convolution3D_CP_2151_elements(319)); -- 
    rr_3677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => type_cast_1577_inst_req_0); -- 
    cr_3682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => type_cast_1577_inst_req_1); -- 
    req_3708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => array_obj_ref_1606_index_offset_req_0); -- 
    req_3713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => array_obj_ref_1606_index_offset_req_1); -- 
    req_3728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => addr_of_1607_final_reg_req_1); -- 
    cr_3778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(319), ack => ptr_deref_1610_store_0_req_1); -- 
    -- CP-element group 320:  merge  fork  transition  place  output  bypass 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	178 
    -- CP-element group 320: 	199 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	200 
    -- CP-element group 320: 	201 
    -- CP-element group 320: 	202 
    -- CP-element group 320:  members (16) 
      -- CP-element group 320: 	 branch_block_stmt_720/merge_stmt_1614_PhiAck/dummy
      -- CP-element group 320: 	 branch_block_stmt_720/merge_stmt_1614__exit__
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626__entry__
      -- CP-element group 320: 	 branch_block_stmt_720/merge_stmt_1614_PhiAck/$exit
      -- CP-element group 320: 	 branch_block_stmt_720/merge_stmt_1614_PhiReqMerge
      -- CP-element group 320: 	 branch_block_stmt_720/merge_stmt_1614_PhiAck/$entry
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/$entry
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_update_start_
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Sample/crr
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Update/$entry
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/call_stmt_1617_Update/ccr
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_sample_start_
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Sample/$entry
      -- CP-element group 320: 	 branch_block_stmt_720/call_stmt_1617_to_assign_stmt_1626/WPIPE_output_pipe_1618_Sample/req
      -- 
    crr_3790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(320), ack => call_stmt_1617_call_req_0); -- 
    ccr_3795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(320), ack => call_stmt_1617_call_req_1); -- 
    req_3804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(320), ack => WPIPE_output_pipe_1618_inst_req_0); -- 
    convolution3D_CP_2151_elements(320) <= OrReduce(convolution3D_CP_2151_elements(178) & convolution3D_CP_2151_elements(199));
    -- CP-element group 321:  transition  output  delay-element  bypass 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	213 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	325 
    -- CP-element group 321:  members (5) 
      -- CP-element group 321: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/$exit
      -- CP-element group 321: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/$exit
      -- CP-element group 321: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/$exit
      -- CP-element group 321: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1678_konst_delay_trans
      -- CP-element group 321: 	 branch_block_stmt_720/ifx_xend_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_req
      -- 
    phi_stmt_1672_req_4623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1672_req_4623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(321), ack => phi_stmt_1672_req_1); -- 
    -- Element group convolution3D_CP_2151_elements(321) is a control-delay.
    cp_element_321_delay: control_delay_element  generic map(name => " 321_delay", delay_value => 1)  port map(req => convolution3D_CP_2151_elements(213), ack => convolution3D_CP_2151_elements(321), clk => clk, reset =>reset);
    -- CP-element group 322:  transition  input  bypass 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	224 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (2) 
      -- CP-element group 322: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Sample/ra
      -- CP-element group 322: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Sample/$exit
      -- 
    ra_4643_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 322_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_0, ack => convolution3D_CP_2151_elements(322)); -- 
    -- CP-element group 323:  transition  input  bypass 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	224 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	324 
    -- CP-element group 323:  members (2) 
      -- CP-element group 323: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Update/ca
      -- CP-element group 323: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/Update/$exit
      -- 
    ca_4648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1675_inst_ack_1, ack => convolution3D_CP_2151_elements(323)); -- 
    -- CP-element group 324:  join  transition  output  bypass 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	323 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	325 
    -- CP-element group 324:  members (6) 
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_req
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/SplitProtocol/$exit
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/type_cast_1675/$exit
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/phi_stmt_1672_sources/$exit
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/phi_stmt_1672/$exit
      -- CP-element group 324: 	 branch_block_stmt_720/whilex_xbody_whilex_xbody_PhiReq/$exit
      -- 
    phi_stmt_1672_req_4649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1672_req_4649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(324), ack => phi_stmt_1672_req_0); -- 
    convolution3D_cp_element_group_324: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convolution3D_cp_element_group_324"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolution3D_CP_2151_elements(322) & convolution3D_CP_2151_elements(323);
      gj_convolution3D_cp_element_group_324 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolution3D_CP_2151_elements(324), clk => clk, reset => reset); --
    end block;
    -- CP-element group 325:  merge  transition  place  bypass 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	321 
    -- CP-element group 325: 	324 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	326 
    -- CP-element group 325:  members (2) 
      -- CP-element group 325: 	 branch_block_stmt_720/merge_stmt_1671_PhiReqMerge
      -- CP-element group 325: 	 branch_block_stmt_720/merge_stmt_1671_PhiAck/$entry
      -- 
    convolution3D_CP_2151_elements(325) <= OrReduce(convolution3D_CP_2151_elements(321) & convolution3D_CP_2151_elements(324));
    -- CP-element group 326:  fork  transition  place  input  output  bypass 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	325 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	220 
    -- CP-element group 326: 	221 
    -- CP-element group 326: 	214 
    -- CP-element group 326: 	218 
    -- CP-element group 326: 	219 
    -- CP-element group 326:  members (20) 
      -- CP-element group 326: 	 branch_block_stmt_720/merge_stmt_1671__exit__
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708__entry__
      -- CP-element group 326: 	 branch_block_stmt_720/merge_stmt_1671_PhiAck/phi_stmt_1672_ack
      -- CP-element group 326: 	 branch_block_stmt_720/merge_stmt_1671_PhiAck/$exit
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/WPIPE_num_out_pipe_1685_Sample/req
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_update_start_
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Sample/crr
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1693_Update/ccr
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_sample_start_
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_update_start_
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Sample/crr
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_720/assign_stmt_1684_to_assign_stmt_1708/call_stmt_1697_Update/ccr
      -- 
    phi_stmt_1672_ack_4654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 326_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1672_ack_0, ack => convolution3D_CP_2151_elements(326)); -- 
    req_3880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(326), ack => WPIPE_num_out_pipe_1685_inst_req_0); -- 
    crr_3908_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3908_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(326), ack => call_stmt_1693_call_req_0); -- 
    ccr_3913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(326), ack => call_stmt_1693_call_req_1); -- 
    crr_3922_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3922_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(326), ack => call_stmt_1697_call_req_0); -- 
    ccr_3927_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3927_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolution3D_CP_2151_elements(326), ack => call_stmt_1697_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar373_1294_resized : std_logic_vector(13 downto 0);
    signal R_indvar373_1294_scaled : std_logic_vector(13 downto 0);
    signal R_indvar379_1010_resized : std_logic_vector(13 downto 0);
    signal R_indvar379_1010_scaled : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1605_resized : std_logic_vector(13 downto 0);
    signal R_ix_x1x_xlcssa_1605_scaled : std_logic_vector(13 downto 0);
    signal add100_1056 : std_logic_vector(63 downto 0);
    signal add106_1074 : std_logic_vector(63 downto 0);
    signal add112_1092 : std_logic_vector(63 downto 0);
    signal add118_1110 : std_logic_vector(63 downto 0);
    signal add124_1128 : std_logic_vector(63 downto 0);
    signal add130_1146 : std_logic_vector(63 downto 0);
    signal add13_770 : std_logic_vector(15 downto 0);
    signal add159_1322 : std_logic_vector(63 downto 0);
    signal add165_1340 : std_logic_vector(63 downto 0);
    signal add171_1358 : std_logic_vector(63 downto 0);
    signal add177_1376 : std_logic_vector(63 downto 0);
    signal add183_1394 : std_logic_vector(63 downto 0);
    signal add189_1412 : std_logic_vector(63 downto 0);
    signal add195_1430 : std_logic_vector(63 downto 0);
    signal add23_795 : std_logic_vector(15 downto 0);
    signal add33_820 : std_logic_vector(15 downto 0);
    signal add43_845 : std_logic_vector(15 downto 0);
    signal add53_870 : std_logic_vector(15 downto 0);
    signal add63_895 : std_logic_vector(31 downto 0);
    signal add73_920 : std_logic_vector(15 downto 0);
    signal add94_1038 : std_logic_vector(63 downto 0);
    signal add_745 : std_logic_vector(31 downto 0);
    signal addx_xi_1545 : std_logic_vector(63 downto 0);
    signal and_1479 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1011_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1011_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1011_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1011_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1011_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1011_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1295_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1606_root_address : std_logic_vector(13 downto 0);
    signal arrayidx199_1297 : std_logic_vector(31 downto 0);
    signal arrayidx211_1608 : std_logic_vector(31 downto 0);
    signal arrayidx_1013 : std_logic_vector(31 downto 0);
    signal call103_1065 : std_logic_vector(7 downto 0);
    signal call109_1083 : std_logic_vector(7 downto 0);
    signal call115_1101 : std_logic_vector(7 downto 0);
    signal call11_761 : std_logic_vector(7 downto 0);
    signal call121_1119 : std_logic_vector(7 downto 0);
    signal call127_1137 : std_logic_vector(7 downto 0);
    signal call152_1300 : std_logic_vector(7 downto 0);
    signal call156_1313 : std_logic_vector(7 downto 0);
    signal call162_1331 : std_logic_vector(7 downto 0);
    signal call168_1349 : std_logic_vector(7 downto 0);
    signal call16_773 : std_logic_vector(7 downto 0);
    signal call174_1367 : std_logic_vector(7 downto 0);
    signal call180_1385 : std_logic_vector(7 downto 0);
    signal call186_1403 : std_logic_vector(7 downto 0);
    signal call192_1421 : std_logic_vector(7 downto 0);
    signal call213_1617 : std_logic_vector(63 downto 0);
    signal call21_786 : std_logic_vector(7 downto 0);
    signal call257_1724 : std_logic_vector(7 downto 0);
    signal call260_1728 : std_logic_vector(7 downto 0);
    signal call262_1731 : std_logic_vector(63 downto 0);
    signal call26_798 : std_logic_vector(7 downto 0);
    signal call2_736 : std_logic_vector(7 downto 0);
    signal call31_811 : std_logic_vector(7 downto 0);
    signal call36_823 : std_logic_vector(7 downto 0);
    signal call41_836 : std_logic_vector(7 downto 0);
    signal call46_848 : std_logic_vector(7 downto 0);
    signal call51_861 : std_logic_vector(7 downto 0);
    signal call56_873 : std_logic_vector(7 downto 0);
    signal call61_886 : std_logic_vector(7 downto 0);
    signal call66_898 : std_logic_vector(7 downto 0);
    signal call6_748 : std_logic_vector(7 downto 0);
    signal call71_911 : std_logic_vector(7 downto 0);
    signal call87_1016 : std_logic_vector(7 downto 0);
    signal call91_1029 : std_logic_vector(7 downto 0);
    signal call97_1047 : std_logic_vector(7 downto 0);
    signal call_723 : std_logic_vector(7 downto 0);
    signal callx_xi_1536 : std_logic_vector(7 downto 0);
    signal cmp149340_1199 : std_logic_vector(0 downto 0);
    signal cmp343_944 : std_logic_vector(0 downto 0);
    signal conv105_1069 : std_logic_vector(63 downto 0);
    signal conv10x_xi_1578 : std_logic_vector(63 downto 0);
    signal conv111_1087 : std_logic_vector(63 downto 0);
    signal conv117_1105 : std_logic_vector(63 downto 0);
    signal conv123_1123 : std_logic_vector(63 downto 0);
    signal conv129_1141 : std_logic_vector(63 downto 0);
    signal conv12_765 : std_logic_vector(15 downto 0);
    signal conv137_1174 : std_logic_vector(31 downto 0);
    signal conv143_1178 : std_logic_vector(31 downto 0);
    signal conv153_1304 : std_logic_vector(63 downto 0);
    signal conv158_1317 : std_logic_vector(63 downto 0);
    signal conv164_1335 : std_logic_vector(63 downto 0);
    signal conv170_1353 : std_logic_vector(63 downto 0);
    signal conv176_1371 : std_logic_vector(63 downto 0);
    signal conv182_1389 : std_logic_vector(63 downto 0);
    signal conv188_1407 : std_logic_vector(63 downto 0);
    signal conv194_1425 : std_logic_vector(63 downto 0);
    signal conv19_777 : std_logic_vector(15 downto 0);
    signal conv1_727 : std_logic_vector(31 downto 0);
    signal conv214_1721 : std_logic_vector(63 downto 0);
    signal conv22_790 : std_logic_vector(15 downto 0);
    signal conv263_1736 : std_logic_vector(63 downto 0);
    signal conv268_1745 : std_logic_vector(31 downto 0);
    signal conv270_1749 : std_logic_vector(31 downto 0);
    signal conv278_1766 : std_logic_vector(7 downto 0);
    signal conv284_1776 : std_logic_vector(7 downto 0);
    signal conv290_1786 : std_logic_vector(7 downto 0);
    signal conv296_1796 : std_logic_vector(7 downto 0);
    signal conv29_802 : std_logic_vector(15 downto 0);
    signal conv302_1806 : std_logic_vector(7 downto 0);
    signal conv308_1816 : std_logic_vector(7 downto 0);
    signal conv314_1826 : std_logic_vector(7 downto 0);
    signal conv320_1836 : std_logic_vector(7 downto 0);
    signal conv32_815 : std_logic_vector(15 downto 0);
    signal conv39_827 : std_logic_vector(15 downto 0);
    signal conv3_740 : std_logic_vector(31 downto 0);
    signal conv42_840 : std_logic_vector(15 downto 0);
    signal conv49_852 : std_logic_vector(15 downto 0);
    signal conv52_865 : std_logic_vector(15 downto 0);
    signal conv59_877 : std_logic_vector(31 downto 0);
    signal conv5x_xi_1540 : std_logic_vector(63 downto 0);
    signal conv62_890 : std_logic_vector(31 downto 0);
    signal conv69_902 : std_logic_vector(15 downto 0);
    signal conv72_915 : std_logic_vector(15 downto 0);
    signal conv79_924 : std_logic_vector(31 downto 0);
    signal conv81_928 : std_logic_vector(31 downto 0);
    signal conv88_1020 : std_logic_vector(63 downto 0);
    signal conv93_1033 : std_logic_vector(63 downto 0);
    signal conv99_1051 : std_logic_vector(63 downto 0);
    signal conv9_752 : std_logic_vector(15 downto 0);
    signal elementx_x015x_xi_1526 : std_logic_vector(63 downto 0);
    signal exitcond22_1445 : std_logic_vector(0 downto 0);
    signal exitcond23_1161 : std_logic_vector(0 downto 0);
    signal exitcond2_1562 : std_logic_vector(0 downto 0);
    signal exitcond_1708 : std_logic_vector(0 downto 0);
    signal iNsTr_17_983 : std_logic_vector(63 downto 0);
    signal incx_xi_1557 : std_logic_vector(7 downto 0);
    signal indvar373_1283 : std_logic_vector(63 downto 0);
    signal indvar379_999 : std_logic_vector(63 downto 0);
    signal indvar_1672 : std_logic_vector(31 downto 0);
    signal indvarx_xnext374_1440 : std_logic_vector(63 downto 0);
    signal indvarx_xnext380_1156 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1703 : std_logic_vector(31 downto 0);
    signal ix_x1x_xlcssa_1466 : std_logic_vector(63 downto 0);
    signal mul138_1183 : std_logic_vector(31 downto 0);
    signal mul141_1188 : std_logic_vector(31 downto 0);
    signal mul144_1193 : std_logic_vector(31 downto 0);
    signal mul241_1684 : std_logic_vector(31 downto 0);
    signal mul271_1754 : std_logic_vector(31 downto 0);
    signal mul274_1759 : std_logic_vector(31 downto 0);
    signal mul82_938 : std_logic_vector(31 downto 0);
    signal mul_933 : std_logic_vector(31 downto 0);
    signal mulx_xi_1590 : std_logic_vector(63 downto 0);
    signal nx_x016x_xi_1519 : std_logic_vector(7 downto 0);
    signal phitmp392_1463 : std_logic_vector(63 downto 0);
    signal ptr_deref_1148_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1148_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1148_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1148_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1148_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1148_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1432_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1432_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1432_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1432_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1432_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1432_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1610_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1610_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1610_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1610_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1610_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1610_word_offset_0 : std_logic_vector(13 downto 0);
    signal sh_promx_xi_1596 : std_logic_vector(63 downto 0);
    signal shl102_1062 : std_logic_vector(63 downto 0);
    signal shl108_1080 : std_logic_vector(63 downto 0);
    signal shl10_758 : std_logic_vector(15 downto 0);
    signal shl114_1098 : std_logic_vector(63 downto 0);
    signal shl120_1116 : std_logic_vector(63 downto 0);
    signal shl126_1134 : std_logic_vector(63 downto 0);
    signal shl12x_xi_1601 : std_logic_vector(63 downto 0);
    signal shl155_1310 : std_logic_vector(63 downto 0);
    signal shl161_1328 : std_logic_vector(63 downto 0);
    signal shl167_1346 : std_logic_vector(63 downto 0);
    signal shl173_1364 : std_logic_vector(63 downto 0);
    signal shl179_1382 : std_logic_vector(63 downto 0);
    signal shl185_1400 : std_logic_vector(63 downto 0);
    signal shl191_1418 : std_logic_vector(63 downto 0);
    signal shl20_783 : std_logic_vector(15 downto 0);
    signal shl30_808 : std_logic_vector(15 downto 0);
    signal shl40_833 : std_logic_vector(15 downto 0);
    signal shl50_858 : std_logic_vector(15 downto 0);
    signal shl60_883 : std_logic_vector(31 downto 0);
    signal shl70_908 : std_logic_vector(15 downto 0);
    signal shl90_1026 : std_logic_vector(63 downto 0);
    signal shl96_1044 : std_logic_vector(63 downto 0);
    signal shl_733 : std_logic_vector(31 downto 0);
    signal shlx_xi_1551 : std_logic_vector(63 downto 0);
    signal shlx_xix_xlcssa_1570 : std_logic_vector(63 downto 0);
    signal shr220338_1633 : std_logic_vector(15 downto 0);
    signal shr281_1772 : std_logic_vector(63 downto 0);
    signal shr287_1782 : std_logic_vector(63 downto 0);
    signal shr293_1792 : std_logic_vector(63 downto 0);
    signal shr299_1802 : std_logic_vector(63 downto 0);
    signal shr305_1812 : std_logic_vector(63 downto 0);
    signal shr311_1822 : std_logic_vector(63 downto 0);
    signal shr317_1832 : std_logic_vector(63 downto 0);
    signal sub_1741 : std_logic_vector(63 downto 0);
    signal subx_xi_1584 : std_logic_vector(63 downto 0);
    signal tmp10_1222 : std_logic_vector(31 downto 0);
    signal tmp11_1227 : std_logic_vector(31 downto 0);
    signal tmp12_1231 : std_logic_vector(31 downto 0);
    signal tmp13_1236 : std_logic_vector(31 downto 0);
    signal tmp14_1240 : std_logic_vector(31 downto 0);
    signal tmp15_1245 : std_logic_vector(31 downto 0);
    signal tmp16_1251 : std_logic_vector(31 downto 0);
    signal tmp17_1257 : std_logic_vector(0 downto 0);
    signal tmp19_1270 : std_logic_vector(31 downto 0);
    signal tmp1_1516 : std_logic_vector(7 downto 0);
    signal tmp20_1274 : std_logic_vector(63 downto 0);
    signal tmp21_1280 : std_logic_vector(63 downto 0);
    signal tmp347_1497 : std_logic_vector(7 downto 0);
    signal tmp349_1502 : std_logic_vector(7 downto 0);
    signal tmp351_1507 : std_logic_vector(7 downto 0);
    signal tmp354_1639 : std_logic_vector(15 downto 0);
    signal tmp371_1212 : std_logic_vector(31 downto 0);
    signal tmp372_1218 : std_logic_vector(0 downto 0);
    signal tmp382_956 : std_logic_vector(31 downto 0);
    signal tmp384_961 : std_logic_vector(31 downto 0);
    signal tmp385_967 : std_logic_vector(31 downto 0);
    signal tmp385x_xop_979 : std_logic_vector(31 downto 0);
    signal tmp386_973 : std_logic_vector(0 downto 0);
    signal tmp390_996 : std_logic_vector(63 downto 0);
    signal tmp3_1643 : std_logic_vector(31 downto 0);
    signal tmp4_1649 : std_logic_vector(31 downto 0);
    signal tmp5_1655 : std_logic_vector(15 downto 0);
    signal tmp6_1660 : std_logic_vector(15 downto 0);
    signal tmp7_1664 : std_logic_vector(31 downto 0);
    signal tmp8_1669 : std_logic_vector(31 downto 0);
    signal tmp_1512 : std_logic_vector(2 downto 0);
    signal tobool_1485 : std_logic_vector(0 downto 0);
    signal type_cast_1003_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1005_wire : std_logic_vector(63 downto 0);
    signal type_cast_1024_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1042_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1060_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1078_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1096_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1114_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1132_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1154_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1197_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1210_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1216_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1249_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1255_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1262_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1278_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1287_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1289_wire : std_logic_vector(63 downto 0);
    signal type_cast_1308_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1326_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1344_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1362_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1398_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1416_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1438_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1457_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1469_wire : std_logic_vector(63 downto 0);
    signal type_cast_1472_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1477_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1522_wire : std_logic_vector(7 downto 0);
    signal type_cast_1525_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1529_wire : std_logic_vector(63 downto 0);
    signal type_cast_1532_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1555_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1573_wire : std_logic_vector(63 downto 0);
    signal type_cast_1581_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1588_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1594_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1631_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1637_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1647_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1653_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1675_wire : std_logic_vector(31 downto 0);
    signal type_cast_1678_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1701_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1719_wire : std_logic_vector(63 downto 0);
    signal type_cast_1734_wire : std_logic_vector(63 downto 0);
    signal type_cast_1770_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1780_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1790_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1800_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1810_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1820_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1830_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_731_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_756_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_781_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_806_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_856_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_881_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_942_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_965_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_971_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_977_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_987_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_994_wire_constant : std_logic_vector(63 downto 0);
    signal umax18_1264 : std_logic_vector(31 downto 0);
    signal umax_1459 : std_logic_vector(31 downto 0);
    signal xx_xop_989 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1011_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1011_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1011_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1011_resized_base_address <= "00000000000000";
    array_obj_ref_1295_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1295_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1295_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1295_resized_base_address <= "00000000000000";
    array_obj_ref_1606_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1606_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1606_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1606_resized_base_address <= "00000000000000";
    ptr_deref_1148_word_offset_0 <= "00000000000000";
    ptr_deref_1432_word_offset_0 <= "00000000000000";
    ptr_deref_1610_word_offset_0 <= "00000000000000";
    type_cast_1003_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1024_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1042_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1060_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1078_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1096_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1132_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1154_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1197_wire_constant <= "00000000000000000000000000000111";
    type_cast_1210_wire_constant <= "00000000000000000000000000000011";
    type_cast_1216_wire_constant <= "00000000000000000000000000000001";
    type_cast_1249_wire_constant <= "00000000000000000000000000000011";
    type_cast_1255_wire_constant <= "00000000000000000000000000000001";
    type_cast_1262_wire_constant <= "00000000000000000000000000000001";
    type_cast_1268_wire_constant <= "11111111111111111111111111111111";
    type_cast_1278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1287_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1308_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1326_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1344_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1362_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1380_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1398_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1416_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1438_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1457_wire_constant <= "00000000000000000000000000000001";
    type_cast_1472_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1477_wire_constant <= "00000000000000000000000000000111";
    type_cast_1483_wire_constant <= "00000000000000000000000000000000";
    type_cast_1525_wire_constant <= "00000000";
    type_cast_1532_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1549_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1555_wire_constant <= "00000001";
    type_cast_1581_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000111";
    type_cast_1588_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000011";
    type_cast_1594_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1631_wire_constant <= "0000000000000011";
    type_cast_1637_wire_constant <= "1111111111111111";
    type_cast_1647_wire_constant <= "00000000000000000000000000000001";
    type_cast_1653_wire_constant <= "0000000000000011";
    type_cast_1678_wire_constant <= "00000000000000000000000000000000";
    type_cast_1701_wire_constant <= "00000000000000000000000000000001";
    type_cast_1770_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1780_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1790_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1800_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1810_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1820_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1830_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_731_wire_constant <= "00000000000000000000000000001000";
    type_cast_756_wire_constant <= "0000000000001000";
    type_cast_781_wire_constant <= "0000000000001000";
    type_cast_806_wire_constant <= "0000000000001000";
    type_cast_831_wire_constant <= "0000000000001000";
    type_cast_856_wire_constant <= "0000000000001000";
    type_cast_881_wire_constant <= "00000000000000000000000000001000";
    type_cast_906_wire_constant <= "0000000000001000";
    type_cast_942_wire_constant <= "00000000000000000000000000000111";
    type_cast_965_wire_constant <= "00000000000000000000000000000011";
    type_cast_971_wire_constant <= "00000000000000000000000000000001";
    type_cast_977_wire_constant <= "11111111111111111111111111111111";
    type_cast_987_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_994_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1283: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1287_wire_constant & type_cast_1289_wire;
      req <= phi_stmt_1283_req_0 & phi_stmt_1283_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1283",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1283_ack_0,
          idata => idata,
          odata => indvar373_1283,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1283
    phi_stmt_1466: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1469_wire & type_cast_1472_wire_constant;
      req <= phi_stmt_1466_req_0 & phi_stmt_1466_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1466",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1466_ack_0,
          idata => idata,
          odata => ix_x1x_xlcssa_1466,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1466
    phi_stmt_1519: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1522_wire & type_cast_1525_wire_constant;
      req <= phi_stmt_1519_req_0 & phi_stmt_1519_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1519",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1519_ack_0,
          idata => idata,
          odata => nx_x016x_xi_1519,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1519
    phi_stmt_1526: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1529_wire & type_cast_1532_wire_constant;
      req <= phi_stmt_1526_req_0 & phi_stmt_1526_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1526",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1526_ack_0,
          idata => idata,
          odata => elementx_x015x_xi_1526,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1526
    phi_stmt_1570: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_1573_wire;
      req(0) <= phi_stmt_1570_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1570",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1570_ack_0,
          idata => idata,
          odata => shlx_xix_xlcssa_1570,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1570
    phi_stmt_1672: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1675_wire & type_cast_1678_wire_constant;
      req <= phi_stmt_1672_req_0 & phi_stmt_1672_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1672",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1672_ack_0,
          idata => idata,
          odata => indvar_1672,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1672
    phi_stmt_999: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1003_wire_constant & type_cast_1005_wire;
      req <= phi_stmt_999_req_0 & phi_stmt_999_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_999",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_999_ack_0,
          idata => idata,
          odata => indvar379_999,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_999
    -- flow-through select operator MUX_1263_inst
    umax18_1264 <= tmp16_1251 when (tmp17_1257(0) /=  '0') else type_cast_1262_wire_constant;
    -- flow-through select operator MUX_1458_inst
    umax_1459 <= tmp371_1212 when (tmp372_1218(0) /=  '0') else type_cast_1457_wire_constant;
    -- flow-through select operator MUX_995_inst
    tmp390_996 <= xx_xop_989 when (tmp386_973(0) /=  '0') else type_cast_994_wire_constant;
    addr_of_1012_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1012_final_reg_req_0;
      addr_of_1012_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1012_final_reg_req_1;
      addr_of_1012_final_reg_ack_1<= rack(0);
      addr_of_1012_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1012_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1011_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1013,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1296_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1296_final_reg_req_0;
      addr_of_1296_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1296_final_reg_req_1;
      addr_of_1296_final_reg_ack_1<= rack(0);
      addr_of_1296_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1296_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1295_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx199_1297,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1607_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1607_final_reg_req_0;
      addr_of_1607_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1607_final_reg_req_1;
      addr_of_1607_final_reg_ack_1<= rack(0);
      addr_of_1607_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1607_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1606_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx211_1608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1005_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1005_inst_req_0;
      type_cast_1005_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1005_inst_req_1;
      type_cast_1005_inst_ack_1<= rack(0);
      type_cast_1005_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1005_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext380_1156,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1005_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1019_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1019_inst_req_0;
      type_cast_1019_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1019_inst_req_1;
      type_cast_1019_inst_ack_1<= rack(0);
      type_cast_1019_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1019_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call87_1016,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_1020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1032_inst_req_0;
      type_cast_1032_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1032_inst_req_1;
      type_cast_1032_inst_ack_1<= rack(0);
      type_cast_1032_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call91_1029,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv93_1033,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1050_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1050_inst_req_0;
      type_cast_1050_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1050_inst_req_1;
      type_cast_1050_inst_ack_1<= rack(0);
      type_cast_1050_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1050_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call97_1047,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv99_1051,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1068_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1068_inst_req_0;
      type_cast_1068_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1068_inst_req_1;
      type_cast_1068_inst_ack_1<= rack(0);
      type_cast_1068_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1068_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call103_1065,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv105_1069,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1086_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1086_inst_req_0;
      type_cast_1086_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1086_inst_req_1;
      type_cast_1086_inst_ack_1<= rack(0);
      type_cast_1086_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1086_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call109_1083,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv111_1087,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1104_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1104_inst_req_0;
      type_cast_1104_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1104_inst_req_1;
      type_cast_1104_inst_ack_1<= rack(0);
      type_cast_1104_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1104_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call115_1101,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv117_1105,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1122_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1122_inst_req_0;
      type_cast_1122_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1122_inst_req_1;
      type_cast_1122_inst_ack_1<= rack(0);
      type_cast_1122_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1122_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call121_1119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv123_1123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1140_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1140_inst_req_0;
      type_cast_1140_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1140_inst_req_1;
      type_cast_1140_inst_ack_1<= rack(0);
      type_cast_1140_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1140_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call127_1137,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv129_1141,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1173_inst_req_0;
      type_cast_1173_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1173_inst_req_1;
      type_cast_1173_inst_ack_1<= rack(0);
      type_cast_1173_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv137_1174,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1177_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1177_inst_req_0;
      type_cast_1177_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1177_inst_req_1;
      type_cast_1177_inst_ack_1<= rack(0);
      type_cast_1177_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1177_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_870,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv143_1178,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1221_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1221_inst_req_0;
      type_cast_1221_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1221_inst_req_1;
      type_cast_1221_inst_ack_1<= rack(0);
      type_cast_1221_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1221_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add53_870,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp10_1222,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1230_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1230_inst_req_0;
      type_cast_1230_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1230_inst_req_1;
      type_cast_1230_inst_ack_1<= rack(0);
      type_cast_1230_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1230_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp12_1231,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1239_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1239_inst_req_0;
      type_cast_1239_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1239_inst_req_1;
      type_cast_1239_inst_ack_1<= rack(0);
      type_cast_1239_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1239_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add73_920,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp14_1240,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1273_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1273_inst_req_0;
      type_cast_1273_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1273_inst_req_1;
      type_cast_1273_inst_ack_1<= rack(0);
      type_cast_1273_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1273_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp19_1270,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp20_1274,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1289_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1289_inst_req_0;
      type_cast_1289_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1289_inst_req_1;
      type_cast_1289_inst_ack_1<= rack(0);
      type_cast_1289_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1289_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext374_1440,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1289_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1303_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1303_inst_req_0;
      type_cast_1303_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1303_inst_req_1;
      type_cast_1303_inst_ack_1<= rack(0);
      type_cast_1303_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1303_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call152_1300,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_1304,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1316_inst_req_0;
      type_cast_1316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1316_inst_req_1;
      type_cast_1316_inst_ack_1<= rack(0);
      type_cast_1316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1316_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call156_1313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv158_1317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1334_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1334_inst_req_0;
      type_cast_1334_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1334_inst_req_1;
      type_cast_1334_inst_ack_1<= rack(0);
      type_cast_1334_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1334_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call162_1331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv164_1335,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1352_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1352_inst_req_0;
      type_cast_1352_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1352_inst_req_1;
      type_cast_1352_inst_ack_1<= rack(0);
      type_cast_1352_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1352_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call168_1349,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv170_1353,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1370_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1370_inst_req_0;
      type_cast_1370_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1370_inst_req_1;
      type_cast_1370_inst_ack_1<= rack(0);
      type_cast_1370_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1370_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call174_1367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv176_1371,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1388_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1388_inst_req_0;
      type_cast_1388_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1388_inst_req_1;
      type_cast_1388_inst_ack_1<= rack(0);
      type_cast_1388_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1388_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call180_1385,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv182_1389,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1406_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1406_inst_req_0;
      type_cast_1406_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1406_inst_req_1;
      type_cast_1406_inst_ack_1<= rack(0);
      type_cast_1406_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1406_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call186_1403,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv188_1407,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1424_inst_req_0;
      type_cast_1424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1424_inst_req_1;
      type_cast_1424_inst_ack_1<= rack(0);
      type_cast_1424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call192_1421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv194_1425,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1462_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1462_inst_req_0;
      type_cast_1462_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1462_inst_req_1;
      type_cast_1462_inst_ack_1<= rack(0);
      type_cast_1462_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1462_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => umax_1459,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => phitmp392_1463,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1469_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1469_inst_req_0;
      type_cast_1469_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1469_inst_req_1;
      type_cast_1469_inst_ack_1<= rack(0);
      type_cast_1469_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1469_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => phitmp392_1463,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1469_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1511_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1511_inst_req_0;
      type_cast_1511_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1511_inst_req_1;
      type_cast_1511_inst_ack_1<= rack(0);
      type_cast_1511_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1511_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp351_1507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp_1512,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1515_inst_req_0;
      type_cast_1515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1515_inst_req_1;
      type_cast_1515_inst_ack_1<= rack(0);
      type_cast_1515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_1512,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp1_1516,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1522_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1522_inst_req_0;
      type_cast_1522_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1522_inst_req_1;
      type_cast_1522_inst_ack_1<= rack(0);
      type_cast_1522_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1522_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => incx_xi_1557,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1522_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1529_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1529_inst_req_0;
      type_cast_1529_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1529_inst_req_1;
      type_cast_1529_inst_ack_1<= rack(0);
      type_cast_1529_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1529_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1529_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1539_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1539_inst_req_0;
      type_cast_1539_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1539_inst_req_1;
      type_cast_1539_inst_ack_1<= rack(0);
      type_cast_1539_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1539_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => callx_xi_1536,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv5x_xi_1540,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1573_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1573_inst_req_0;
      type_cast_1573_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1573_inst_req_1;
      type_cast_1573_inst_ack_1<= rack(0);
      type_cast_1573_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1573_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shlx_xi_1551,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1573_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1577_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1577_inst_req_0;
      type_cast_1577_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1577_inst_req_1;
      type_cast_1577_inst_ack_1<= rack(0);
      type_cast_1577_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1577_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul144_1193,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10x_xi_1578,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1642_inst_req_0;
      type_cast_1642_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1642_inst_req_1;
      type_cast_1642_inst_ack_1<= rack(0);
      type_cast_1642_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1642_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp354_1639,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp3_1643,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1663_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1663_inst_req_0;
      type_cast_1663_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1663_inst_req_1;
      type_cast_1663_inst_ack_1<= rack(0);
      type_cast_1663_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1663_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_1660,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_1664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1675_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1675_inst_req_0;
      type_cast_1675_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1675_inst_req_1;
      type_cast_1675_inst_ack_1<= rack(0);
      type_cast_1675_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1675_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1703,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1675_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1720_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1720_inst_req_0;
      type_cast_1720_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1720_inst_req_1;
      type_cast_1720_inst_ack_1<= rack(0);
      type_cast_1720_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1720_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1719_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv214_1721,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1735_inst_req_0;
      type_cast_1735_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1735_inst_req_1;
      type_cast_1735_inst_ack_1<= rack(0);
      type_cast_1735_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1735_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1734_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv263_1736,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1744_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1744_inst_req_0;
      type_cast_1744_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1744_inst_req_1;
      type_cast_1744_inst_ack_1<= rack(0);
      type_cast_1744_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1744_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add43_845,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv268_1745,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1748_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1748_inst_req_0;
      type_cast_1748_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1748_inst_req_1;
      type_cast_1748_inst_ack_1<= rack(0);
      type_cast_1748_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1748_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add33_820,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv270_1749,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1765_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1765_inst_req_0;
      type_cast_1765_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1765_inst_req_1;
      type_cast_1765_inst_ack_1<= rack(0);
      type_cast_1765_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1765_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => sub_1741,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv278_1766,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1775_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1775_inst_req_0;
      type_cast_1775_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1775_inst_req_1;
      type_cast_1775_inst_ack_1<= rack(0);
      type_cast_1775_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1775_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr281_1772,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv284_1776,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1785_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1785_inst_req_0;
      type_cast_1785_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1785_inst_req_1;
      type_cast_1785_inst_ack_1<= rack(0);
      type_cast_1785_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1785_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr287_1782,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv290_1786,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1795_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1795_inst_req_0;
      type_cast_1795_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1795_inst_req_1;
      type_cast_1795_inst_ack_1<= rack(0);
      type_cast_1795_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1795_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr293_1792,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv296_1796,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1805_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1805_inst_req_0;
      type_cast_1805_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1805_inst_req_1;
      type_cast_1805_inst_ack_1<= rack(0);
      type_cast_1805_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1805_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr299_1802,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv302_1806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1815_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1815_inst_req_0;
      type_cast_1815_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1815_inst_req_1;
      type_cast_1815_inst_ack_1<= rack(0);
      type_cast_1815_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1815_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr305_1812,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv308_1816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1825_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1825_inst_req_0;
      type_cast_1825_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1825_inst_req_1;
      type_cast_1825_inst_ack_1<= rack(0);
      type_cast_1825_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1825_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr311_1822,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv314_1826,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1835_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1835_inst_req_0;
      type_cast_1835_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1835_inst_req_1;
      type_cast_1835_inst_ack_1<= rack(0);
      type_cast_1835_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1835_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr317_1832,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv320_1836,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_726_inst_req_0;
      type_cast_726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_726_inst_req_1;
      type_cast_726_inst_ack_1<= rack(0);
      type_cast_726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_723,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv1_727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_739_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_739_inst_req_0;
      type_cast_739_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_739_inst_req_1;
      type_cast_739_inst_ack_1<= rack(0);
      type_cast_739_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_739_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call2_736,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_751_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_751_inst_req_1;
      type_cast_751_inst_ack_1<= rack(0);
      type_cast_751_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_751_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call6_748,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9_752,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_764_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_764_inst_req_0;
      type_cast_764_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_764_inst_req_1;
      type_cast_764_inst_ack_1<= rack(0);
      type_cast_764_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_764_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call11_761,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_765,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_776_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_776_inst_req_0;
      type_cast_776_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_776_inst_req_1;
      type_cast_776_inst_ack_1<= rack(0);
      type_cast_776_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_776_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call16_773,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_777,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_789_inst_req_0;
      type_cast_789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_789_inst_req_1;
      type_cast_789_inst_ack_1<= rack(0);
      type_cast_789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call21_786,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_801_inst_req_0;
      type_cast_801_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_801_inst_req_1;
      type_cast_801_inst_ack_1<= rack(0);
      type_cast_801_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_801_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call26_798,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_802,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_814_inst_req_0;
      type_cast_814_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_814_inst_req_1;
      type_cast_814_inst_ack_1<= rack(0);
      type_cast_814_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_814_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call31_811,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv32_815,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_826_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_826_inst_req_0;
      type_cast_826_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_826_inst_req_1;
      type_cast_826_inst_ack_1<= rack(0);
      type_cast_826_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_826_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call36_823,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv39_827,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_839_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_839_inst_req_0;
      type_cast_839_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_839_inst_req_1;
      type_cast_839_inst_ack_1<= rack(0);
      type_cast_839_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_839_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call41_836,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_840,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_851_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_851_inst_req_0;
      type_cast_851_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_851_inst_req_1;
      type_cast_851_inst_ack_1<= rack(0);
      type_cast_851_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_851_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call46_848,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv49_852,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_864_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_864_inst_req_0;
      type_cast_864_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_864_inst_req_1;
      type_cast_864_inst_ack_1<= rack(0);
      type_cast_864_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_864_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call51_861,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv52_865,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_876_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_876_inst_req_0;
      type_cast_876_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_876_inst_req_1;
      type_cast_876_inst_ack_1<= rack(0);
      type_cast_876_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_876_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call56_873,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv59_877,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_889_inst_req_0;
      type_cast_889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_889_inst_req_1;
      type_cast_889_inst_ack_1<= rack(0);
      type_cast_889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call61_886,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv62_890,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_901_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_901_inst_req_0;
      type_cast_901_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_901_inst_req_1;
      type_cast_901_inst_ack_1<= rack(0);
      type_cast_901_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_901_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call66_898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_902,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_914_inst_req_0;
      type_cast_914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_914_inst_req_1;
      type_cast_914_inst_ack_1<= rack(0);
      type_cast_914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call71_911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv72_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_923_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_923_inst_req_1;
      type_cast_923_inst_ack_1<= rack(0);
      type_cast_923_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_923_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add13_770,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_924,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_927_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_927_inst_req_0;
      type_cast_927_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_927_inst_req_1;
      type_cast_927_inst_ack_1<= rack(0);
      type_cast_927_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_927_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => add23_795,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv81_928,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_982_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_982_inst_req_0;
      type_cast_982_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_982_inst_req_1;
      type_cast_982_inst_ack_1<= rack(0);
      type_cast_982_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_982_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp385x_xop_979,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_17_983,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1011_index_1_rename
    process(R_indvar379_1010_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar379_1010_resized;
      ov(13 downto 0) := iv;
      R_indvar379_1010_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1011_index_1_resize
    process(indvar379_999) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar379_999;
      ov := iv(13 downto 0);
      R_indvar379_1010_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1011_root_address_inst
    process(array_obj_ref_1011_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1011_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1011_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1295_index_1_rename
    process(R_indvar373_1294_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar373_1294_resized;
      ov(13 downto 0) := iv;
      R_indvar373_1294_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1295_index_1_resize
    process(indvar373_1283) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar373_1283;
      ov := iv(13 downto 0);
      R_indvar373_1294_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1295_root_address_inst
    process(array_obj_ref_1295_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1295_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1295_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1606_index_1_rename
    process(R_ix_x1x_xlcssa_1605_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_ix_x1x_xlcssa_1605_resized;
      ov(13 downto 0) := iv;
      R_ix_x1x_xlcssa_1605_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1606_index_1_resize
    process(ix_x1x_xlcssa_1466) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ix_x1x_xlcssa_1466;
      ov := iv(13 downto 0);
      R_ix_x1x_xlcssa_1605_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1606_root_address_inst
    process(array_obj_ref_1606_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1606_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1606_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1148_addr_0
    process(ptr_deref_1148_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1148_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1148_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1148_base_resize
    process(arrayidx_1013) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1013;
      ov := iv(13 downto 0);
      ptr_deref_1148_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1148_gather_scatter
    process(add130_1146) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add130_1146;
      ov(63 downto 0) := iv;
      ptr_deref_1148_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1148_root_address_inst
    process(ptr_deref_1148_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1148_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1148_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_addr_0
    process(ptr_deref_1432_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1432_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1432_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_base_resize
    process(arrayidx199_1297) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx199_1297;
      ov := iv(13 downto 0);
      ptr_deref_1432_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_gather_scatter
    process(add195_1430) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add195_1430;
      ov(63 downto 0) := iv;
      ptr_deref_1432_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1432_root_address_inst
    process(ptr_deref_1432_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1432_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1432_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1610_addr_0
    process(ptr_deref_1610_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1610_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1610_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1610_base_resize
    process(arrayidx211_1608) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx211_1608;
      ov := iv(13 downto 0);
      ptr_deref_1610_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1610_gather_scatter
    process(shl12x_xi_1601) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := shl12x_xi_1601;
      ov(63 downto 0) := iv;
      ptr_deref_1610_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1610_root_address_inst
    process(ptr_deref_1610_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1610_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1610_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1162_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond23_1161;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1162_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1162_branch_req_0,
          ack0 => if_stmt_1162_branch_ack_0,
          ack1 => if_stmt_1162_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1200_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp149340_1199;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1200_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1200_branch_req_0,
          ack0 => if_stmt_1200_branch_ack_0,
          ack1 => if_stmt_1200_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1446_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond22_1445;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1446_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1446_branch_req_0,
          ack0 => if_stmt_1446_branch_ack_0,
          ack1 => if_stmt_1446_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1486_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tobool_1485;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1486_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1486_branch_req_0,
          ack0 => if_stmt_1486_branch_ack_0,
          ack1 => if_stmt_1486_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1563_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond2_1562;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1563_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1563_branch_req_0,
          ack0 => if_stmt_1563_branch_ack_0,
          ack1 => if_stmt_1563_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1709_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1708;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1709_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1709_branch_req_0,
          ack0 => if_stmt_1709_branch_ack_0,
          ack1 => if_stmt_1709_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_945_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp343_944;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_945_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_945_branch_req_0,
          ack0 => if_stmt_945_branch_ack_0,
          ack1 => if_stmt_945_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1638_inst
    process(add53_870) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(add53_870, type_cast_1637_wire_constant, tmp_var);
      tmp354_1639 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1269_inst
    process(umax18_1264) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(umax18_1264, type_cast_1268_wire_constant, tmp_var);
      tmp19_1270 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1648_inst
    process(tmp3_1643) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp3_1643, type_cast_1647_wire_constant, tmp_var);
      tmp4_1649 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1702_inst
    process(indvar_1672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1672, type_cast_1701_wire_constant, tmp_var);
      indvarx_xnext_1703 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_978_inst
    process(tmp385_967) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp385_967, type_cast_977_wire_constant, tmp_var);
      tmp385x_xop_979 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1155_inst
    process(indvar379_999) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar379_999, type_cast_1154_wire_constant, tmp_var);
      indvarx_xnext380_1156 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1279_inst
    process(tmp20_1274) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp20_1274, type_cast_1278_wire_constant, tmp_var);
      tmp21_1280 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1439_inst
    process(indvar373_1283) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar373_1283, type_cast_1438_wire_constant, tmp_var);
      indvarx_xnext374_1440 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_988_inst
    process(iNsTr_17_983) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_17_983, type_cast_987_wire_constant, tmp_var);
      xx_xop_989 <= tmp_var; --
    end process;
    -- binary operator ADD_u8_u8_1556_inst
    process(nx_x016x_xi_1519) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(nx_x016x_xi_1519, type_cast_1555_wire_constant, tmp_var);
      incx_xi_1557 <= tmp_var; --
    end process;
    -- binary operator AND_u32_u32_1478_inst
    process(mul144_1193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mul144_1193, type_cast_1477_wire_constant, tmp_var);
      and_1479 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_1595_inst
    process(mulx_xi_1590) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(mulx_xi_1590, type_cast_1594_wire_constant, tmp_var);
      sh_promx_xi_1596 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1484_inst
    process(and_1479) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(and_1479, type_cast_1483_wire_constant, tmp_var);
      tobool_1485 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1707_inst
    process(indvarx_xnext_1703, tmp4_1649) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1703, tmp4_1649, tmp_var);
      exitcond_1708 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1160_inst
    process(indvarx_xnext380_1156, tmp390_996) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext380_1156, tmp390_996, tmp_var);
      exitcond23_1161 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1444_inst
    process(indvarx_xnext374_1440, tmp21_1280) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext374_1440, tmp21_1280, tmp_var);
      exitcond22_1445 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1561_inst
    process(incx_xi_1557, tmp1_1516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(incx_xi_1557, tmp1_1516, tmp_var);
      exitcond2_1562 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1632_inst
    process(add23_795) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add23_795, type_cast_1631_wire_constant, tmp_var);
      shr220338_1633 <= tmp_var; --
    end process;
    -- binary operator LSHR_u16_u16_1654_inst
    process(add23_795) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(add23_795, type_cast_1653_wire_constant, tmp_var);
      tmp5_1655 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1211_inst
    process(mul144_1193) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul144_1193, type_cast_1210_wire_constant, tmp_var);
      tmp371_1212 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1250_inst
    process(tmp15_1245) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp15_1245, type_cast_1249_wire_constant, tmp_var);
      tmp16_1251 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_966_inst
    process(tmp384_961) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp384_961, type_cast_965_wire_constant, tmp_var);
      tmp385_967 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1771_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1770_wire_constant, tmp_var);
      shr281_1772 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1781_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1780_wire_constant, tmp_var);
      shr287_1782 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1791_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1790_wire_constant, tmp_var);
      shr293_1792 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1801_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1800_wire_constant, tmp_var);
      shr299_1802 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1811_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1810_wire_constant, tmp_var);
      shr305_1812 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1821_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1820_wire_constant, tmp_var);
      shr311_1822 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1831_inst
    process(sub_1741) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(sub_1741, type_cast_1830_wire_constant, tmp_var);
      shr317_1832 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1659_inst
    process(add73_920, tmp5_1655) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(add73_920, tmp5_1655, tmp_var);
      tmp6_1660 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1182_inst
    process(conv143_1178, conv81_928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv143_1178, conv81_928, tmp_var);
      mul138_1183 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1187_inst
    process(mul138_1183, add63_895) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul138_1183, add63_895, tmp_var);
      mul141_1188 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1192_inst
    process(mul141_1188, conv137_1174) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul141_1188, conv137_1174, tmp_var);
      mul144_1193 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1226_inst
    process(add63_895, tmp10_1222) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_895, tmp10_1222, tmp_var);
      tmp11_1227 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1235_inst
    process(tmp11_1227, tmp12_1231) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp11_1227, tmp12_1231, tmp_var);
      tmp13_1236 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1244_inst
    process(tmp13_1236, tmp14_1240) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_1236, tmp14_1240, tmp_var);
      tmp15_1245 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1668_inst
    process(add63_895, tmp7_1664) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add63_895, tmp7_1664, tmp_var);
      tmp8_1669 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1683_inst
    process(tmp8_1669, indvar_1672) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp8_1669, indvar_1672, tmp_var);
      mul241_1684 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1753_inst
    process(conv268_1745, conv270_1749) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv268_1745, conv270_1749, tmp_var);
      mul271_1754 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1758_inst
    process(mul271_1754, conv143_1178) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul271_1754, conv143_1178, tmp_var);
      mul274_1759 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_932_inst
    process(conv79_924, add_745) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv79_924, add_745, tmp_var);
      mul_933 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_937_inst
    process(mul_933, conv81_928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_933, conv81_928, tmp_var);
      mul82_938 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_955_inst
    process(add_745, conv79_924) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_745, conv79_924, tmp_var);
      tmp382_956 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_960_inst
    process(tmp382_956, conv81_928) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp382_956, conv81_928, tmp_var);
      tmp384_961 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_1496_inst
    process(call51_861, call21_786) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(call51_861, call21_786, tmp_var);
      tmp347_1497 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_1501_inst
    process(tmp347_1497, call61_886) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp347_1497, call61_886, tmp_var);
      tmp349_1502 <= tmp_var; --
    end process;
    -- binary operator MUL_u8_u8_1506_inst
    process(tmp349_1502, call71_911) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp349_1502, call71_911, tmp_var);
      tmp351_1507 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_769_inst
    process(shl10_758, conv12_765) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl10_758, conv12_765, tmp_var);
      add13_770 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_794_inst
    process(shl20_783, conv22_790) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl20_783, conv22_790, tmp_var);
      add23_795 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_819_inst
    process(shl30_808, conv32_815) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl30_808, conv32_815, tmp_var);
      add33_820 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_844_inst
    process(shl40_833, conv42_840) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl40_833, conv42_840, tmp_var);
      add43_845 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_869_inst
    process(shl50_858, conv52_865) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl50_858, conv52_865, tmp_var);
      add53_870 <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_919_inst
    process(shl70_908, conv72_915) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl70_908, conv72_915, tmp_var);
      add73_920 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_744_inst
    process(shl_733, conv3_740) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_733, conv3_740, tmp_var);
      add_745 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_894_inst
    process(shl60_883, conv62_890) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl60_883, conv62_890, tmp_var);
      add63_895 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1037_inst
    process(shl90_1026, conv93_1033) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl90_1026, conv93_1033, tmp_var);
      add94_1038 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1055_inst
    process(shl96_1044, conv99_1051) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl96_1044, conv99_1051, tmp_var);
      add100_1056 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1073_inst
    process(shl102_1062, conv105_1069) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl102_1062, conv105_1069, tmp_var);
      add106_1074 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1091_inst
    process(shl108_1080, conv111_1087) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl108_1080, conv111_1087, tmp_var);
      add112_1092 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1109_inst
    process(shl114_1098, conv117_1105) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl114_1098, conv117_1105, tmp_var);
      add118_1110 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1127_inst
    process(shl120_1116, conv123_1123) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl120_1116, conv123_1123, tmp_var);
      add124_1128 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1145_inst
    process(shl126_1134, conv129_1141) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl126_1134, conv129_1141, tmp_var);
      add130_1146 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1321_inst
    process(shl155_1310, conv158_1317) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl155_1310, conv158_1317, tmp_var);
      add159_1322 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1339_inst
    process(shl161_1328, conv164_1335) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl161_1328, conv164_1335, tmp_var);
      add165_1340 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1357_inst
    process(shl167_1346, conv170_1353) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl167_1346, conv170_1353, tmp_var);
      add171_1358 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1375_inst
    process(shl173_1364, conv176_1371) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl173_1364, conv176_1371, tmp_var);
      add177_1376 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1393_inst
    process(shl179_1382, conv182_1389) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl179_1382, conv182_1389, tmp_var);
      add183_1394 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1411_inst
    process(shl185_1400, conv188_1407) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl185_1400, conv188_1407, tmp_var);
      add189_1412 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1429_inst
    process(shl191_1418, conv194_1425) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl191_1418, conv194_1425, tmp_var);
      add195_1430 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_1544_inst
    process(conv5x_xi_1540, elementx_x015x_xi_1526) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(conv5x_xi_1540, elementx_x015x_xi_1526, tmp_var);
      addx_xi_1545 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_757_inst
    process(conv9_752) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv9_752, type_cast_756_wire_constant, tmp_var);
      shl10_758 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_782_inst
    process(conv19_777) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv19_777, type_cast_781_wire_constant, tmp_var);
      shl20_783 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_807_inst
    process(conv29_802) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv29_802, type_cast_806_wire_constant, tmp_var);
      shl30_808 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_832_inst
    process(conv39_827) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv39_827, type_cast_831_wire_constant, tmp_var);
      shl40_833 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_857_inst
    process(conv49_852) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv49_852, type_cast_856_wire_constant, tmp_var);
      shl50_858 <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_907_inst
    process(conv69_902) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv69_902, type_cast_906_wire_constant, tmp_var);
      shl70_908 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_732_inst
    process(conv1_727) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv1_727, type_cast_731_wire_constant, tmp_var);
      shl_733 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_882_inst
    process(conv59_877) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv59_877, type_cast_881_wire_constant, tmp_var);
      shl60_883 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1025_inst
    process(conv88_1020) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv88_1020, type_cast_1024_wire_constant, tmp_var);
      shl90_1026 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1043_inst
    process(add94_1038) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add94_1038, type_cast_1042_wire_constant, tmp_var);
      shl96_1044 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1061_inst
    process(add100_1056) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add100_1056, type_cast_1060_wire_constant, tmp_var);
      shl102_1062 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1079_inst
    process(add106_1074) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add106_1074, type_cast_1078_wire_constant, tmp_var);
      shl108_1080 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1097_inst
    process(add112_1092) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add112_1092, type_cast_1096_wire_constant, tmp_var);
      shl114_1098 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1115_inst
    process(add118_1110) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add118_1110, type_cast_1114_wire_constant, tmp_var);
      shl120_1116 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1133_inst
    process(add124_1128) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add124_1128, type_cast_1132_wire_constant, tmp_var);
      shl126_1134 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1309_inst
    process(conv153_1304) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv153_1304, type_cast_1308_wire_constant, tmp_var);
      shl155_1310 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1327_inst
    process(add159_1322) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add159_1322, type_cast_1326_wire_constant, tmp_var);
      shl161_1328 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1345_inst
    process(add165_1340) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add165_1340, type_cast_1344_wire_constant, tmp_var);
      shl167_1346 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1363_inst
    process(add171_1358) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add171_1358, type_cast_1362_wire_constant, tmp_var);
      shl173_1364 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1381_inst
    process(add177_1376) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add177_1376, type_cast_1380_wire_constant, tmp_var);
      shl179_1382 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1399_inst
    process(add183_1394) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add183_1394, type_cast_1398_wire_constant, tmp_var);
      shl185_1400 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1417_inst
    process(add189_1412) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add189_1412, type_cast_1416_wire_constant, tmp_var);
      shl191_1418 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1550_inst
    process(addx_xi_1545) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(addx_xi_1545, type_cast_1549_wire_constant, tmp_var);
      shlx_xi_1551 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1589_inst
    process(subx_xi_1584) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(subx_xi_1584, type_cast_1588_wire_constant, tmp_var);
      mulx_xi_1590 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_1600_inst
    process(shlx_xix_xlcssa_1570, sh_promx_xi_1596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(shlx_xix_xlcssa_1570, sh_promx_xi_1596, tmp_var);
      shl12x_xi_1601 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1583_inst
    process(type_cast_1581_wire_constant, conv10x_xi_1578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(type_cast_1581_wire_constant, conv10x_xi_1578, tmp_var);
      subx_xi_1584 <= tmp_var; --
    end process;
    -- binary operator SUB_u64_u64_1740_inst
    process(conv263_1736, conv214_1721) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSub_proc(conv263_1736, conv214_1721, tmp_var);
      sub_1741 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1198_inst
    process(mul144_1193) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul144_1193, type_cast_1197_wire_constant, tmp_var);
      cmp149340_1199 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1217_inst
    process(tmp371_1212) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp371_1212, type_cast_1216_wire_constant, tmp_var);
      tmp372_1218 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1256_inst
    process(tmp16_1251) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp16_1251, type_cast_1255_wire_constant, tmp_var);
      tmp17_1257 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_943_inst
    process(mul82_938) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul82_938, type_cast_942_wire_constant, tmp_var);
      cmp343_944 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_972_inst
    process(tmp385_967) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp385_967, type_cast_971_wire_constant, tmp_var);
      tmp386_973 <= tmp_var; --
    end process;
    -- shared split operator group (102) : array_obj_ref_1011_index_offset 
    ApIntAdd_group_102: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar379_1010_scaled;
      array_obj_ref_1011_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1011_index_offset_req_0;
      array_obj_ref_1011_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1011_index_offset_req_1;
      array_obj_ref_1011_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_102_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_102_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_102",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 102
    -- shared split operator group (103) : array_obj_ref_1295_index_offset 
    ApIntAdd_group_103: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar373_1294_scaled;
      array_obj_ref_1295_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1295_index_offset_req_0;
      array_obj_ref_1295_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1295_index_offset_req_1;
      array_obj_ref_1295_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_103_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_103_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_103",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 103
    -- shared split operator group (104) : array_obj_ref_1606_index_offset 
    ApIntAdd_group_104: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_ix_x1x_xlcssa_1605_scaled;
      array_obj_ref_1606_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1606_index_offset_req_0;
      array_obj_ref_1606_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1606_index_offset_req_1;
      array_obj_ref_1606_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_104_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_104_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_104",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 104
    -- unary operator type_cast_1719_inst
    process(call213_1617) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call213_1617, tmp_var);
      type_cast_1719_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1734_inst
    process(call262_1731) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", call262_1731, tmp_var);
      type_cast_1734_wire <= tmp_var; -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1148_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1148_store_0_req_0;
      ptr_deref_1148_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1148_store_0_req_1;
      ptr_deref_1148_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1148_word_address_0;
      data_in <= ptr_deref_1148_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(13 downto 0),
          mdata => memory_space_2_sr_data(63 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1432_store_0 ptr_deref_1610_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1432_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1610_store_0_req_0;
      ptr_deref_1432_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1610_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1432_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1610_store_0_req_1;
      ptr_deref_1432_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1610_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup1_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup1_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1432_word_address_0 & ptr_deref_1610_word_address_0;
      data_in <= ptr_deref_1432_data_0 & ptr_deref_1610_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(13 downto 0),
          mdata => memory_space_1_sr_data(63 downto 0),
          mtag => memory_space_1_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : RPIPE_input_done_pipe_1723_inst RPIPE_input_done_pipe_1727_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_input_done_pipe_1723_inst_req_0;
      reqL_unguarded(0) <= RPIPE_input_done_pipe_1727_inst_req_0;
      RPIPE_input_done_pipe_1723_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_input_done_pipe_1727_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_input_done_pipe_1723_inst_req_1;
      reqR_unguarded(0) <= RPIPE_input_done_pipe_1727_inst_req_1;
      RPIPE_input_done_pipe_1723_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_input_done_pipe_1727_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      call257_1724 <= data_out(15 downto 8);
      call260_1728 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_maxpool_input_pipe_847_inst RPIPE_maxpool_input_pipe_860_inst RPIPE_maxpool_input_pipe_810_inst RPIPE_maxpool_input_pipe_872_inst RPIPE_maxpool_input_pipe_910_inst RPIPE_maxpool_input_pipe_885_inst RPIPE_maxpool_input_pipe_722_inst RPIPE_maxpool_input_pipe_835_inst RPIPE_maxpool_input_pipe_897_inst RPIPE_maxpool_input_pipe_735_inst RPIPE_maxpool_input_pipe_785_inst RPIPE_maxpool_input_pipe_822_inst RPIPE_maxpool_input_pipe_797_inst RPIPE_maxpool_input_pipe_1046_inst RPIPE_maxpool_input_pipe_1384_inst RPIPE_maxpool_input_pipe_1366_inst RPIPE_maxpool_input_pipe_1348_inst RPIPE_maxpool_input_pipe_1330_inst RPIPE_maxpool_input_pipe_1312_inst RPIPE_maxpool_input_pipe_1299_inst RPIPE_maxpool_input_pipe_772_inst RPIPE_maxpool_input_pipe_1015_inst RPIPE_maxpool_input_pipe_1028_inst RPIPE_maxpool_input_pipe_1420_inst RPIPE_maxpool_input_pipe_760_inst RPIPE_maxpool_input_pipe_1402_inst RPIPE_maxpool_input_pipe_1136_inst RPIPE_maxpool_input_pipe_1118_inst RPIPE_maxpool_input_pipe_1100_inst RPIPE_maxpool_input_pipe_1082_inst RPIPE_maxpool_input_pipe_747_inst RPIPE_maxpool_input_pipe_1064_inst RPIPE_maxpool_input_pipe_1535_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(263 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 32 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 32 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 32 downto 0);
      signal guard_vector : std_logic_vector( 32 downto 0);
      constant outBUFs : IntegerArray(32 downto 0) := (32 => 1, 31 => 1, 30 => 1, 29 => 1, 28 => 1, 27 => 1, 26 => 1, 25 => 1, 24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(32 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false, 25 => false, 26 => false, 27 => false, 28 => false, 29 => false, 30 => false, 31 => false, 32 => false);
      constant guardBuffering: IntegerArray(32 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2, 25 => 2, 26 => 2, 27 => 2, 28 => 2, 29 => 2, 30 => 2, 31 => 2, 32 => 2);
      -- 
    begin -- 
      reqL_unguarded(32) <= RPIPE_maxpool_input_pipe_847_inst_req_0;
      reqL_unguarded(31) <= RPIPE_maxpool_input_pipe_860_inst_req_0;
      reqL_unguarded(30) <= RPIPE_maxpool_input_pipe_810_inst_req_0;
      reqL_unguarded(29) <= RPIPE_maxpool_input_pipe_872_inst_req_0;
      reqL_unguarded(28) <= RPIPE_maxpool_input_pipe_910_inst_req_0;
      reqL_unguarded(27) <= RPIPE_maxpool_input_pipe_885_inst_req_0;
      reqL_unguarded(26) <= RPIPE_maxpool_input_pipe_722_inst_req_0;
      reqL_unguarded(25) <= RPIPE_maxpool_input_pipe_835_inst_req_0;
      reqL_unguarded(24) <= RPIPE_maxpool_input_pipe_897_inst_req_0;
      reqL_unguarded(23) <= RPIPE_maxpool_input_pipe_735_inst_req_0;
      reqL_unguarded(22) <= RPIPE_maxpool_input_pipe_785_inst_req_0;
      reqL_unguarded(21) <= RPIPE_maxpool_input_pipe_822_inst_req_0;
      reqL_unguarded(20) <= RPIPE_maxpool_input_pipe_797_inst_req_0;
      reqL_unguarded(19) <= RPIPE_maxpool_input_pipe_1046_inst_req_0;
      reqL_unguarded(18) <= RPIPE_maxpool_input_pipe_1384_inst_req_0;
      reqL_unguarded(17) <= RPIPE_maxpool_input_pipe_1366_inst_req_0;
      reqL_unguarded(16) <= RPIPE_maxpool_input_pipe_1348_inst_req_0;
      reqL_unguarded(15) <= RPIPE_maxpool_input_pipe_1330_inst_req_0;
      reqL_unguarded(14) <= RPIPE_maxpool_input_pipe_1312_inst_req_0;
      reqL_unguarded(13) <= RPIPE_maxpool_input_pipe_1299_inst_req_0;
      reqL_unguarded(12) <= RPIPE_maxpool_input_pipe_772_inst_req_0;
      reqL_unguarded(11) <= RPIPE_maxpool_input_pipe_1015_inst_req_0;
      reqL_unguarded(10) <= RPIPE_maxpool_input_pipe_1028_inst_req_0;
      reqL_unguarded(9) <= RPIPE_maxpool_input_pipe_1420_inst_req_0;
      reqL_unguarded(8) <= RPIPE_maxpool_input_pipe_760_inst_req_0;
      reqL_unguarded(7) <= RPIPE_maxpool_input_pipe_1402_inst_req_0;
      reqL_unguarded(6) <= RPIPE_maxpool_input_pipe_1136_inst_req_0;
      reqL_unguarded(5) <= RPIPE_maxpool_input_pipe_1118_inst_req_0;
      reqL_unguarded(4) <= RPIPE_maxpool_input_pipe_1100_inst_req_0;
      reqL_unguarded(3) <= RPIPE_maxpool_input_pipe_1082_inst_req_0;
      reqL_unguarded(2) <= RPIPE_maxpool_input_pipe_747_inst_req_0;
      reqL_unguarded(1) <= RPIPE_maxpool_input_pipe_1064_inst_req_0;
      reqL_unguarded(0) <= RPIPE_maxpool_input_pipe_1535_inst_req_0;
      RPIPE_maxpool_input_pipe_847_inst_ack_0 <= ackL_unguarded(32);
      RPIPE_maxpool_input_pipe_860_inst_ack_0 <= ackL_unguarded(31);
      RPIPE_maxpool_input_pipe_810_inst_ack_0 <= ackL_unguarded(30);
      RPIPE_maxpool_input_pipe_872_inst_ack_0 <= ackL_unguarded(29);
      RPIPE_maxpool_input_pipe_910_inst_ack_0 <= ackL_unguarded(28);
      RPIPE_maxpool_input_pipe_885_inst_ack_0 <= ackL_unguarded(27);
      RPIPE_maxpool_input_pipe_722_inst_ack_0 <= ackL_unguarded(26);
      RPIPE_maxpool_input_pipe_835_inst_ack_0 <= ackL_unguarded(25);
      RPIPE_maxpool_input_pipe_897_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_maxpool_input_pipe_735_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_maxpool_input_pipe_785_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_maxpool_input_pipe_822_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_maxpool_input_pipe_797_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_maxpool_input_pipe_1046_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_maxpool_input_pipe_1384_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_maxpool_input_pipe_1366_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_maxpool_input_pipe_1348_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_maxpool_input_pipe_1330_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_maxpool_input_pipe_1312_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_maxpool_input_pipe_1299_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_maxpool_input_pipe_772_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_maxpool_input_pipe_1015_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_maxpool_input_pipe_1028_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_maxpool_input_pipe_1420_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_maxpool_input_pipe_760_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_maxpool_input_pipe_1402_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_maxpool_input_pipe_1136_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_maxpool_input_pipe_1118_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_maxpool_input_pipe_1100_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_maxpool_input_pipe_1082_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_maxpool_input_pipe_747_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_maxpool_input_pipe_1064_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_maxpool_input_pipe_1535_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(32) <= RPIPE_maxpool_input_pipe_847_inst_req_1;
      reqR_unguarded(31) <= RPIPE_maxpool_input_pipe_860_inst_req_1;
      reqR_unguarded(30) <= RPIPE_maxpool_input_pipe_810_inst_req_1;
      reqR_unguarded(29) <= RPIPE_maxpool_input_pipe_872_inst_req_1;
      reqR_unguarded(28) <= RPIPE_maxpool_input_pipe_910_inst_req_1;
      reqR_unguarded(27) <= RPIPE_maxpool_input_pipe_885_inst_req_1;
      reqR_unguarded(26) <= RPIPE_maxpool_input_pipe_722_inst_req_1;
      reqR_unguarded(25) <= RPIPE_maxpool_input_pipe_835_inst_req_1;
      reqR_unguarded(24) <= RPIPE_maxpool_input_pipe_897_inst_req_1;
      reqR_unguarded(23) <= RPIPE_maxpool_input_pipe_735_inst_req_1;
      reqR_unguarded(22) <= RPIPE_maxpool_input_pipe_785_inst_req_1;
      reqR_unguarded(21) <= RPIPE_maxpool_input_pipe_822_inst_req_1;
      reqR_unguarded(20) <= RPIPE_maxpool_input_pipe_797_inst_req_1;
      reqR_unguarded(19) <= RPIPE_maxpool_input_pipe_1046_inst_req_1;
      reqR_unguarded(18) <= RPIPE_maxpool_input_pipe_1384_inst_req_1;
      reqR_unguarded(17) <= RPIPE_maxpool_input_pipe_1366_inst_req_1;
      reqR_unguarded(16) <= RPIPE_maxpool_input_pipe_1348_inst_req_1;
      reqR_unguarded(15) <= RPIPE_maxpool_input_pipe_1330_inst_req_1;
      reqR_unguarded(14) <= RPIPE_maxpool_input_pipe_1312_inst_req_1;
      reqR_unguarded(13) <= RPIPE_maxpool_input_pipe_1299_inst_req_1;
      reqR_unguarded(12) <= RPIPE_maxpool_input_pipe_772_inst_req_1;
      reqR_unguarded(11) <= RPIPE_maxpool_input_pipe_1015_inst_req_1;
      reqR_unguarded(10) <= RPIPE_maxpool_input_pipe_1028_inst_req_1;
      reqR_unguarded(9) <= RPIPE_maxpool_input_pipe_1420_inst_req_1;
      reqR_unguarded(8) <= RPIPE_maxpool_input_pipe_760_inst_req_1;
      reqR_unguarded(7) <= RPIPE_maxpool_input_pipe_1402_inst_req_1;
      reqR_unguarded(6) <= RPIPE_maxpool_input_pipe_1136_inst_req_1;
      reqR_unguarded(5) <= RPIPE_maxpool_input_pipe_1118_inst_req_1;
      reqR_unguarded(4) <= RPIPE_maxpool_input_pipe_1100_inst_req_1;
      reqR_unguarded(3) <= RPIPE_maxpool_input_pipe_1082_inst_req_1;
      reqR_unguarded(2) <= RPIPE_maxpool_input_pipe_747_inst_req_1;
      reqR_unguarded(1) <= RPIPE_maxpool_input_pipe_1064_inst_req_1;
      reqR_unguarded(0) <= RPIPE_maxpool_input_pipe_1535_inst_req_1;
      RPIPE_maxpool_input_pipe_847_inst_ack_1 <= ackR_unguarded(32);
      RPIPE_maxpool_input_pipe_860_inst_ack_1 <= ackR_unguarded(31);
      RPIPE_maxpool_input_pipe_810_inst_ack_1 <= ackR_unguarded(30);
      RPIPE_maxpool_input_pipe_872_inst_ack_1 <= ackR_unguarded(29);
      RPIPE_maxpool_input_pipe_910_inst_ack_1 <= ackR_unguarded(28);
      RPIPE_maxpool_input_pipe_885_inst_ack_1 <= ackR_unguarded(27);
      RPIPE_maxpool_input_pipe_722_inst_ack_1 <= ackR_unguarded(26);
      RPIPE_maxpool_input_pipe_835_inst_ack_1 <= ackR_unguarded(25);
      RPIPE_maxpool_input_pipe_897_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_maxpool_input_pipe_735_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_maxpool_input_pipe_785_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_maxpool_input_pipe_822_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_maxpool_input_pipe_797_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_maxpool_input_pipe_1046_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_maxpool_input_pipe_1384_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_maxpool_input_pipe_1366_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_maxpool_input_pipe_1348_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_maxpool_input_pipe_1330_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_maxpool_input_pipe_1312_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_maxpool_input_pipe_1299_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_maxpool_input_pipe_772_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_maxpool_input_pipe_1015_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_maxpool_input_pipe_1028_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_maxpool_input_pipe_1420_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_maxpool_input_pipe_760_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_maxpool_input_pipe_1402_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_maxpool_input_pipe_1136_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_maxpool_input_pipe_1118_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_maxpool_input_pipe_1100_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_maxpool_input_pipe_1082_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_maxpool_input_pipe_747_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_maxpool_input_pipe_1064_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_maxpool_input_pipe_1535_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      guard_vector(25)  <=  '1';
      guard_vector(26)  <=  '1';
      guard_vector(27)  <=  '1';
      guard_vector(28)  <=  '1';
      guard_vector(29)  <=  '1';
      guard_vector(30)  <=  '1';
      guard_vector(31)  <=  '1';
      guard_vector(32)  <=  '1';
      call46_848 <= data_out(263 downto 256);
      call51_861 <= data_out(255 downto 248);
      call31_811 <= data_out(247 downto 240);
      call56_873 <= data_out(239 downto 232);
      call71_911 <= data_out(231 downto 224);
      call61_886 <= data_out(223 downto 216);
      call_723 <= data_out(215 downto 208);
      call41_836 <= data_out(207 downto 200);
      call66_898 <= data_out(199 downto 192);
      call2_736 <= data_out(191 downto 184);
      call21_786 <= data_out(183 downto 176);
      call36_823 <= data_out(175 downto 168);
      call26_798 <= data_out(167 downto 160);
      call97_1047 <= data_out(159 downto 152);
      call180_1385 <= data_out(151 downto 144);
      call174_1367 <= data_out(143 downto 136);
      call168_1349 <= data_out(135 downto 128);
      call162_1331 <= data_out(127 downto 120);
      call156_1313 <= data_out(119 downto 112);
      call152_1300 <= data_out(111 downto 104);
      call16_773 <= data_out(103 downto 96);
      call87_1016 <= data_out(95 downto 88);
      call91_1029 <= data_out(87 downto 80);
      call192_1421 <= data_out(79 downto 72);
      call11_761 <= data_out(71 downto 64);
      call186_1403 <= data_out(63 downto 56);
      call127_1137 <= data_out(55 downto 48);
      call121_1119 <= data_out(47 downto 40);
      call115_1101 <= data_out(39 downto 32);
      call109_1083 <= data_out(31 downto 24);
      call6_748 <= data_out(23 downto 16);
      call103_1065 <= data_out(15 downto 8);
      callx_xi_1536 <= data_out(7 downto 0);
      maxpool_input_pipe_read_1_gI: SplitGuardInterface generic map(name => "maxpool_input_pipe_read_1_gI", nreqs => 33, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      maxpool_input_pipe_read_1: InputPortRevised -- 
        generic map ( name => "maxpool_input_pipe_read_1", data_width => 8,  num_reqs => 33,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => maxpool_input_pipe_pipe_read_req(0),
          oack => maxpool_input_pipe_pipe_read_ack(0),
          odata => maxpool_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_1837_inst WPIPE_maxpool_output_pipe_1840_inst WPIPE_maxpool_output_pipe_1843_inst WPIPE_maxpool_output_pipe_1846_inst WPIPE_maxpool_output_pipe_1849_inst WPIPE_maxpool_output_pipe_1852_inst WPIPE_maxpool_output_pipe_1855_inst WPIPE_maxpool_output_pipe_1858_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1837_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1840_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1843_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1846_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1849_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1852_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1855_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1858_inst_req_0;
      WPIPE_maxpool_output_pipe_1837_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1840_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1843_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1846_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1849_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1852_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1855_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1858_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_1837_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_1840_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_1843_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_1846_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_1849_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_1852_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_1855_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_1858_inst_req_1;
      WPIPE_maxpool_output_pipe_1837_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_1840_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_1843_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_1846_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_1849_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_1852_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_1855_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_1858_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv320_1836 & conv314_1826 & conv308_1816 & conv302_1806 & conv296_1796 & conv290_1786 & conv284_1776 & conv278_1766;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_num_out_pipe_1685_inst WPIPE_num_out_pipe_1688_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_num_out_pipe_1685_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_num_out_pipe_1688_inst_req_0;
      WPIPE_num_out_pipe_1685_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_num_out_pipe_1688_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_num_out_pipe_1685_inst_req_1;
      update_req_unguarded(0) <= WPIPE_num_out_pipe_1688_inst_req_1;
      WPIPE_num_out_pipe_1685_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_num_out_pipe_1688_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= add33_820 & add43_845;
      num_out_pipe_write_1_gI: SplitGuardInterface generic map(name => "num_out_pipe_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "num_out_pipe", data_width => 16, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => num_out_pipe_pipe_write_req(0),
          oack => num_out_pipe_pipe_write_ack(0),
          odata => num_out_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_output_pipe_1618_inst WPIPE_output_pipe_1621_inst WPIPE_output_pipe_1624_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal sample_req, sample_ack : BooleanArray( 2 downto 0);
      signal update_req, update_ack : BooleanArray( 2 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 2 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      sample_req_unguarded(2) <= WPIPE_output_pipe_1618_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_output_pipe_1621_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_output_pipe_1624_inst_req_0;
      WPIPE_output_pipe_1618_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_output_pipe_1621_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_output_pipe_1624_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(2) <= WPIPE_output_pipe_1618_inst_req_1;
      update_req_unguarded(1) <= WPIPE_output_pipe_1621_inst_req_1;
      update_req_unguarded(0) <= WPIPE_output_pipe_1624_inst_req_1;
      WPIPE_output_pipe_1618_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_output_pipe_1621_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_output_pipe_1624_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      data_in <= add33_820 & add43_845 & add53_870;
      output_pipe_write_2_gI: SplitGuardInterface generic map(name => "output_pipe_write_2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_2: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 3, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared call operator group (0) : call_stmt_1617_call call_stmt_1731_call 
    timer_call_group_0: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1617_call_req_0;
      reqL_unguarded(0) <= call_stmt_1731_call_req_0;
      call_stmt_1617_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1731_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1617_call_req_1;
      reqR_unguarded(0) <= call_stmt_1731_call_req_1;
      call_stmt_1617_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1731_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      timer_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      timer_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "timer_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      timer_call_group_0_gI: SplitGuardInterface generic map(name => "timer_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call213_1617 <= data_out(127 downto 64);
      call262_1731 <= data_out(63 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 2,
        nreqs => 2,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => timer_call_reqs(0),
          ackR => timer_call_acks(0),
          tagR => timer_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => timer_return_acks(0), -- cross-over
          ackL => timer_return_reqs(0), -- cross-over
          dataL => timer_return_data(63 downto 0),
          tagL => timer_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1693_call 
    loadKernelChannel_call_group_1: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1693_call_req_0;
      call_stmt_1693_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1693_call_req_1;
      call_stmt_1693_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadKernelChannel_call_group_1_gI: SplitGuardInterface generic map(name => "loadKernelChannel_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul241_1684 & shr220338_1633;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadKernelChannel_call_reqs(0),
          ackR => loadKernelChannel_call_acks(0),
          dataR => loadKernelChannel_call_data(47 downto 0),
          tagR => loadKernelChannel_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => loadKernelChannel_return_acks(0), -- cross-over
          ackL => loadKernelChannel_return_reqs(0), -- cross-over
          tagL => loadKernelChannel_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1697_call 
    access_T_call_group_2: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1697_call_req_0;
      call_stmt_1697_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1697_call_req_1;
      call_stmt_1697_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      access_T_call_group_2_gI: SplitGuardInterface generic map(name => "access_T_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= add33_820 & shr220338_1633 & add13_770;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 48,
        owidth => 48,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => access_T_call_reqs(0),
          ackR => access_T_call_acks(0),
          dataR => access_T_call_data(47 downto 0),
          tagR => access_T_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => access_T_return_acks(0), -- cross-over
          ackL => access_T_return_reqs(0), -- cross-over
          tagL => access_T_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1761_call 
    sendB_call_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1761_call_req_0;
      call_stmt_1761_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1761_call_req_1;
      call_stmt_1761_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendB_call_group_3_gI: SplitGuardInterface generic map(name => "sendB_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= mul274_1759;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => sendB_call_reqs(0),
          ackR => sendB_call_acks(0),
          dataR => sendB_call_data(31 downto 0),
          tagR => sendB_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendB_return_acks(0), -- cross-over
          ackL => sendB_return_reqs(0), -- cross-over
          tagL => sendB_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end convolution3D_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convolve is -- 
  generic (tag_length : integer); 
  port ( -- 
    input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe2_pipe_read_data : in   std_logic_vector(63 downto 0);
    input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe3_pipe_read_data : in   std_logic_vector(63 downto 0);
    input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe1_pipe_read_data : in   std_logic_vector(63 downto 0);
    kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_read_data : in   std_logic_vector(63 downto 0);
    kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_read_data : in   std_logic_vector(63 downto 0);
    input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_pipe4_pipe_read_data : in   std_logic_vector(63 downto 0);
    kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_read_data : in   std_logic_vector(63 downto 0);
    num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convolve;
architecture convolve_arch of convolve is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convolve_CP_4675_start: Boolean;
  signal convolve_CP_4675_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal slice_2105_inst_req_0 : boolean;
  signal slice_2097_inst_req_0 : boolean;
  signal slice_2117_inst_req_1 : boolean;
  signal slice_2129_inst_ack_0 : boolean;
  signal slice_2089_inst_req_0 : boolean;
  signal n_col_3054_1912_buf_ack_0 : boolean;
  signal nacc2_3080_1902_buf_ack_0 : boolean;
  signal phi_stmt_1913_req_0 : boolean;
  signal slice_2097_inst_ack_0 : boolean;
  signal slice_2105_inst_ack_1 : boolean;
  signal slice_2125_inst_req_1 : boolean;
  signal slice_2093_inst_ack_0 : boolean;
  signal nacc2_3080_1902_buf_req_0 : boolean;
  signal slice_2089_inst_ack_0 : boolean;
  signal slice_2105_inst_req_1 : boolean;
  signal slice_2093_inst_req_0 : boolean;
  signal phi_stmt_1908_ack_0 : boolean;
  signal n_chl_3032_1923_buf_ack_0 : boolean;
  signal phi_stmt_1903_req_1 : boolean;
  signal phi_stmt_1919_req_0 : boolean;
  signal phi_stmt_1913_req_1 : boolean;
  signal n_num_3043_1918_buf_ack_0 : boolean;
  signal phi_stmt_1919_ack_0 : boolean;
  signal n_row_3062_1907_buf_req_0 : boolean;
  signal phi_stmt_1903_req_0 : boolean;
  signal n_row_3062_1907_buf_ack_0 : boolean;
  signal n_col_3054_1912_buf_req_1 : boolean;
  signal phi_stmt_1919_req_1 : boolean;
  signal n_row_3062_1907_buf_req_1 : boolean;
  signal n_col_3054_1912_buf_ack_1 : boolean;
  signal n_row_3062_1907_buf_ack_1 : boolean;
  signal phi_stmt_1908_req_1 : boolean;
  signal n_chl_3032_1923_buf_req_0 : boolean;
  signal nacc2_3080_1902_buf_req_1 : boolean;
  signal phi_stmt_1913_ack_0 : boolean;
  signal n_num_3043_1918_buf_req_0 : boolean;
  signal n_num_3043_1918_buf_req_1 : boolean;
  signal nacc2_3080_1902_buf_ack_1 : boolean;
  signal phi_stmt_1903_ack_0 : boolean;
  signal n_num_3043_1918_buf_ack_1 : boolean;
  signal phi_stmt_1908_req_0 : boolean;
  signal n_col_3054_1912_buf_req_0 : boolean;
  signal slice_2113_inst_req_0 : boolean;
  signal slice_2105_inst_ack_0 : boolean;
  signal slice_2121_inst_req_0 : boolean;
  signal slice_2113_inst_ack_0 : boolean;
  signal slice_2097_inst_req_1 : boolean;
  signal slice_2113_inst_ack_1 : boolean;
  signal slice_2121_inst_ack_0 : boolean;
  signal slice_2125_inst_ack_1 : boolean;
  signal slice_2097_inst_ack_1 : boolean;
  signal slice_2109_inst_req_0 : boolean;
  signal slice_2089_inst_req_1 : boolean;
  signal slice_2129_inst_req_1 : boolean;
  signal slice_2101_inst_req_0 : boolean;
  signal slice_2101_inst_ack_0 : boolean;
  signal slice_2093_inst_req_1 : boolean;
  signal slice_2093_inst_ack_1 : boolean;
  signal slice_2109_inst_ack_0 : boolean;
  signal slice_2089_inst_ack_1 : boolean;
  signal slice_2113_inst_req_1 : boolean;
  signal slice_2117_inst_ack_1 : boolean;
  signal slice_2117_inst_req_0 : boolean;
  signal slice_2125_inst_req_0 : boolean;
  signal slice_2125_inst_ack_0 : boolean;
  signal slice_2129_inst_ack_1 : boolean;
  signal slice_2129_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1876_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1876_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1876_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1876_inst_ack_1 : boolean;
  signal SUB_u16_u16_1878_inst_req_0 : boolean;
  signal SUB_u16_u16_1878_inst_ack_0 : boolean;
  signal SUB_u16_u16_1878_inst_req_1 : boolean;
  signal SUB_u16_u16_1878_inst_ack_1 : boolean;
  signal RPIPE_num_out_pipe_1881_inst_req_0 : boolean;
  signal RPIPE_num_out_pipe_1881_inst_ack_0 : boolean;
  signal RPIPE_num_out_pipe_1881_inst_req_1 : boolean;
  signal RPIPE_num_out_pipe_1881_inst_ack_1 : boolean;
  signal SUB_u16_u16_1883_inst_req_0 : boolean;
  signal SUB_u16_u16_1883_inst_ack_0 : boolean;
  signal SUB_u16_u16_1883_inst_req_1 : boolean;
  signal SUB_u16_u16_1883_inst_ack_1 : boolean;
  signal RPIPE_size_pipe_1886_inst_req_0 : boolean;
  signal RPIPE_size_pipe_1886_inst_ack_0 : boolean;
  signal RPIPE_size_pipe_1886_inst_req_1 : boolean;
  signal RPIPE_size_pipe_1886_inst_ack_1 : boolean;
  signal SUB_u16_u16_1888_inst_req_0 : boolean;
  signal SUB_u16_u16_1888_inst_ack_0 : boolean;
  signal SUB_u16_u16_1888_inst_req_1 : boolean;
  signal SUB_u16_u16_1888_inst_ack_1 : boolean;
  signal do_while_stmt_1890_branch_req_0 : boolean;
  signal phi_stmt_1892_req_1 : boolean;
  signal phi_stmt_1892_req_0 : boolean;
  signal phi_stmt_1892_ack_0 : boolean;
  signal nacc1_3071_1897_buf_req_0 : boolean;
  signal nacc1_3071_1897_buf_ack_0 : boolean;
  signal nacc1_3071_1897_buf_req_1 : boolean;
  signal nacc1_3071_1897_buf_ack_1 : boolean;
  signal phi_stmt_1898_req_1 : boolean;
  signal phi_stmt_1898_req_0 : boolean;
  signal phi_stmt_1898_ack_0 : boolean;
  signal n_chl_3032_1923_buf_req_1 : boolean;
  signal n_chl_3032_1923_buf_ack_1 : boolean;
  signal RPIPE_input_pipe1_1936_inst_req_0 : boolean;
  signal RPIPE_input_pipe1_1936_inst_ack_0 : boolean;
  signal RPIPE_input_pipe1_1936_inst_req_1 : boolean;
  signal RPIPE_input_pipe1_1936_inst_ack_1 : boolean;
  signal RPIPE_input_pipe2_1940_inst_req_0 : boolean;
  signal RPIPE_input_pipe2_1940_inst_ack_0 : boolean;
  signal RPIPE_input_pipe2_1940_inst_req_1 : boolean;
  signal RPIPE_input_pipe2_1940_inst_ack_1 : boolean;
  signal RPIPE_input_pipe3_1944_inst_req_0 : boolean;
  signal RPIPE_input_pipe3_1944_inst_ack_0 : boolean;
  signal RPIPE_input_pipe3_1944_inst_req_1 : boolean;
  signal RPIPE_input_pipe3_1944_inst_ack_1 : boolean;
  signal RPIPE_input_pipe4_1948_inst_req_0 : boolean;
  signal RPIPE_input_pipe4_1948_inst_ack_0 : boolean;
  signal RPIPE_input_pipe4_1948_inst_req_1 : boolean;
  signal RPIPE_input_pipe4_1948_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1952_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1952_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_1 : boolean;
  signal slice_2101_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1956_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1956_inst_req_1 : boolean;
  signal slice_2109_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_1 : boolean;
  signal slice_2117_inst_ack_0 : boolean;
  signal slice_2121_inst_ack_1 : boolean;
  signal slice_2121_inst_req_1 : boolean;
  signal slice_2101_inst_req_1 : boolean;
  signal slice_2109_inst_req_1 : boolean;
  signal slice_2133_inst_req_0 : boolean;
  signal slice_2133_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1960_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1960_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_1 : boolean;
  signal slice_2437_inst_req_0 : boolean;
  signal slice_2405_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3008_inst_ack_1 : boolean;
  signal slice_2449_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_1964_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_1964_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_1 : boolean;
  signal slice_2425_inst_req_0 : boolean;
  signal SUB_u16_u16_2986_inst_req_1 : boolean;
  signal slice_2405_inst_ack_0 : boolean;
  signal slice_2425_inst_ack_0 : boolean;
  signal W_read_ip_1946_delayed_1_0_1966_inst_req_0 : boolean;
  signal W_read_ip_1946_delayed_1_0_1966_inst_ack_0 : boolean;
  signal W_read_ip_1946_delayed_1_0_1966_inst_req_1 : boolean;
  signal slice_2437_inst_ack_0 : boolean;
  signal W_read_ip_1946_delayed_1_0_1966_inst_ack_1 : boolean;
  signal slice_2397_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3008_inst_ack_0 : boolean;
  signal slice_2397_inst_ack_1 : boolean;
  signal slice_2445_inst_req_0 : boolean;
  signal W_read_ip_1952_delayed_1_0_1975_inst_req_0 : boolean;
  signal W_read_ip_1952_delayed_1_0_1975_inst_ack_0 : boolean;
  signal W_read_ip_1952_delayed_1_0_1975_inst_req_1 : boolean;
  signal W_read_ip_1952_delayed_1_0_1975_inst_ack_1 : boolean;
  signal slice_2445_inst_ack_0 : boolean;
  signal slice_2413_inst_req_0 : boolean;
  signal W_read_ip_1958_delayed_1_0_1984_inst_req_0 : boolean;
  signal W_read_ip_1958_delayed_1_0_1984_inst_ack_0 : boolean;
  signal W_read_ip_1958_delayed_1_0_1984_inst_req_1 : boolean;
  signal W_read_ip_1958_delayed_1_0_1984_inst_ack_1 : boolean;
  signal slice_2425_inst_req_1 : boolean;
  signal slice_2413_inst_ack_0 : boolean;
  signal W_read_ip_1964_delayed_1_0_1993_inst_req_0 : boolean;
  signal W_read_ip_1964_delayed_1_0_1993_inst_ack_0 : boolean;
  signal W_read_ip_1964_delayed_1_0_1993_inst_req_1 : boolean;
  signal slice_2437_inst_req_1 : boolean;
  signal W_read_ip_1964_delayed_1_0_1993_inst_ack_1 : boolean;
  signal slice_2405_inst_req_1 : boolean;
  signal slice_2425_inst_ack_1 : boolean;
  signal W_acc2_2893_delayed_2_0_2949_inst_req_0 : boolean;
  signal W_write_input_1978_delayed_1_0_2011_inst_req_0 : boolean;
  signal slice_2437_inst_ack_1 : boolean;
  signal W_write_input_1978_delayed_1_0_2011_inst_ack_0 : boolean;
  signal W_write_input_1978_delayed_1_0_2011_inst_req_1 : boolean;
  signal W_write_input_1978_delayed_1_0_2011_inst_ack_1 : boolean;
  signal slice_2401_inst_req_0 : boolean;
  signal SUB_u16_u16_2986_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2015_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2015_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3008_inst_req_0 : boolean;
  signal slice_2413_inst_req_1 : boolean;
  signal slice_2413_inst_ack_1 : boolean;
  signal W_acc2_2893_delayed_2_0_2949_inst_ack_0 : boolean;
  signal W_write_input_1982_delayed_1_0_2018_inst_req_0 : boolean;
  signal W_write_input_1982_delayed_1_0_2018_inst_ack_0 : boolean;
  signal W_write_input_1982_delayed_1_0_2018_inst_req_1 : boolean;
  signal W_write_input_1982_delayed_1_0_2018_inst_ack_1 : boolean;
  signal W_store_kernel_2941_delayed_1_0_3004_inst_req_1 : boolean;
  signal slice_2401_inst_ack_0 : boolean;
  signal slice_2445_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2022_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2022_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_1 : boolean;
  signal W_acc1_2884_delayed_2_0_2937_inst_req_0 : boolean;
  signal W_write_input_1986_delayed_1_0_2025_inst_req_0 : boolean;
  signal W_write_input_1986_delayed_1_0_2025_inst_ack_0 : boolean;
  signal W_acc2_2893_delayed_2_0_2949_inst_req_1 : boolean;
  signal W_write_input_1986_delayed_1_0_2025_inst_req_1 : boolean;
  signal W_write_input_1986_delayed_1_0_2025_inst_ack_1 : boolean;
  signal slice_2417_inst_req_0 : boolean;
  signal slice_2441_inst_req_0 : boolean;
  signal W_store_kernel_2941_delayed_1_0_3004_inst_ack_1 : boolean;
  signal slice_2449_inst_req_0 : boolean;
  signal slice_2417_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2029_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_0 : boolean;
  signal slice_2429_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2029_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_1 : boolean;
  signal slice_2429_inst_ack_0 : boolean;
  signal slice_2401_inst_req_1 : boolean;
  signal W_write_input_1990_delayed_1_0_2032_inst_req_0 : boolean;
  signal slice_2441_inst_ack_0 : boolean;
  signal W_write_input_1990_delayed_1_0_2032_inst_ack_0 : boolean;
  signal W_acc2_2893_delayed_2_0_2949_inst_ack_1 : boolean;
  signal W_write_input_1990_delayed_1_0_2032_inst_req_1 : boolean;
  signal W_write_input_1990_delayed_1_0_2032_inst_ack_1 : boolean;
  signal slice_2405_inst_ack_1 : boolean;
  signal W_acc1_2884_delayed_2_0_2937_inst_ack_0 : boolean;
  signal slice_2429_inst_req_1 : boolean;
  signal slice_2417_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2036_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2036_inst_req_1 : boolean;
  signal slice_2441_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_1 : boolean;
  signal W_store_kernel_2941_delayed_1_0_3004_inst_req_0 : boolean;
  signal slice_2417_inst_ack_1 : boolean;
  signal slice_2429_inst_ack_1 : boolean;
  signal W_store_kernel_2941_delayed_1_0_3004_inst_ack_0 : boolean;
  signal slice_2441_inst_ack_1 : boolean;
  signal slice_2445_inst_ack_1 : boolean;
  signal slice_2401_inst_ack_1 : boolean;
  signal slice_2041_inst_req_0 : boolean;
  signal slice_2041_inst_ack_0 : boolean;
  signal slice_2041_inst_req_1 : boolean;
  signal slice_2041_inst_ack_1 : boolean;
  signal slice_2045_inst_req_0 : boolean;
  signal slice_2045_inst_ack_0 : boolean;
  signal slice_2045_inst_req_1 : boolean;
  signal slice_2045_inst_ack_1 : boolean;
  signal slice_2049_inst_req_0 : boolean;
  signal slice_2049_inst_ack_0 : boolean;
  signal slice_2049_inst_req_1 : boolean;
  signal slice_2049_inst_ack_1 : boolean;
  signal slice_2053_inst_req_0 : boolean;
  signal slice_2053_inst_ack_0 : boolean;
  signal slice_2053_inst_req_1 : boolean;
  signal slice_2053_inst_ack_1 : boolean;
  signal slice_2057_inst_req_0 : boolean;
  signal slice_2057_inst_ack_0 : boolean;
  signal slice_2057_inst_req_1 : boolean;
  signal slice_2057_inst_ack_1 : boolean;
  signal slice_2061_inst_req_0 : boolean;
  signal slice_2061_inst_ack_0 : boolean;
  signal slice_2061_inst_req_1 : boolean;
  signal slice_2061_inst_ack_1 : boolean;
  signal slice_2065_inst_req_0 : boolean;
  signal slice_2065_inst_ack_0 : boolean;
  signal slice_2065_inst_req_1 : boolean;
  signal slice_2065_inst_ack_1 : boolean;
  signal slice_2069_inst_req_0 : boolean;
  signal slice_2069_inst_ack_0 : boolean;
  signal slice_2069_inst_req_1 : boolean;
  signal slice_2069_inst_ack_1 : boolean;
  signal slice_2073_inst_req_0 : boolean;
  signal slice_2073_inst_ack_0 : boolean;
  signal slice_2073_inst_req_1 : boolean;
  signal slice_2073_inst_ack_1 : boolean;
  signal slice_2077_inst_req_0 : boolean;
  signal slice_2077_inst_ack_0 : boolean;
  signal slice_2077_inst_req_1 : boolean;
  signal slice_2077_inst_ack_1 : boolean;
  signal slice_2081_inst_req_0 : boolean;
  signal slice_2081_inst_ack_0 : boolean;
  signal slice_2081_inst_req_1 : boolean;
  signal slice_2081_inst_ack_1 : boolean;
  signal slice_2085_inst_req_0 : boolean;
  signal slice_2085_inst_ack_0 : boolean;
  signal slice_2085_inst_req_1 : boolean;
  signal slice_2085_inst_ack_1 : boolean;
  signal slice_2133_inst_req_1 : boolean;
  signal slice_2133_inst_ack_1 : boolean;
  signal slice_2137_inst_req_0 : boolean;
  signal slice_2137_inst_ack_0 : boolean;
  signal slice_2137_inst_req_1 : boolean;
  signal slice_2137_inst_ack_1 : boolean;
  signal slice_2141_inst_req_0 : boolean;
  signal slice_2141_inst_ack_0 : boolean;
  signal slice_2141_inst_req_1 : boolean;
  signal slice_2141_inst_ack_1 : boolean;
  signal slice_2145_inst_req_0 : boolean;
  signal slice_2145_inst_ack_0 : boolean;
  signal slice_2145_inst_req_1 : boolean;
  signal slice_2145_inst_ack_1 : boolean;
  signal slice_2149_inst_req_0 : boolean;
  signal slice_2149_inst_ack_0 : boolean;
  signal slice_2149_inst_req_1 : boolean;
  signal slice_2149_inst_ack_1 : boolean;
  signal slice_2153_inst_req_0 : boolean;
  signal slice_2153_inst_ack_0 : boolean;
  signal slice_2153_inst_req_1 : boolean;
  signal slice_2153_inst_ack_1 : boolean;
  signal slice_2157_inst_req_0 : boolean;
  signal slice_2157_inst_ack_0 : boolean;
  signal slice_2157_inst_req_1 : boolean;
  signal slice_2157_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k1_3008_inst_req_1 : boolean;
  signal slice_2161_inst_req_0 : boolean;
  signal slice_2161_inst_ack_0 : boolean;
  signal W_acc1_2884_delayed_2_0_2937_inst_ack_1 : boolean;
  signal slice_2161_inst_req_1 : boolean;
  signal slice_2161_inst_ack_1 : boolean;
  signal slice_2409_inst_ack_1 : boolean;
  signal slice_2409_inst_req_1 : boolean;
  signal slice_2449_inst_ack_1 : boolean;
  signal slice_2421_inst_ack_1 : boolean;
  signal W_acc1_2884_delayed_2_0_2937_inst_req_1 : boolean;
  signal slice_2165_inst_req_0 : boolean;
  signal slice_2165_inst_ack_0 : boolean;
  signal slice_2165_inst_req_1 : boolean;
  signal slice_2165_inst_ack_1 : boolean;
  signal slice_2409_inst_ack_0 : boolean;
  signal slice_2397_inst_ack_0 : boolean;
  signal slice_2449_inst_req_1 : boolean;
  signal slice_2421_inst_req_1 : boolean;
  signal slice_2409_inst_req_0 : boolean;
  signal slice_2397_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe1_2306_inst_req_0 : boolean;
  signal slice_2433_inst_ack_1 : boolean;
  signal RPIPE_kernel_pipe1_2306_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe1_2306_inst_req_1 : boolean;
  signal slice_2433_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe1_2306_inst_ack_1 : boolean;
  signal SUB_u16_u16_2986_inst_ack_0 : boolean;
  signal SUB_u16_u16_2986_inst_req_0 : boolean;
  signal slice_2421_inst_ack_0 : boolean;
  signal slice_2421_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2310_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe2_2310_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2310_inst_req_1 : boolean;
  signal slice_2433_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe2_2310_inst_ack_1 : boolean;
  signal slice_2433_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_2314_inst_req_0 : boolean;
  signal RPIPE_kernel_pipe3_2314_inst_ack_0 : boolean;
  signal RPIPE_kernel_pipe3_2314_inst_req_1 : boolean;
  signal RPIPE_kernel_pipe3_2314_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2318_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2318_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2318_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k1_2318_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2322_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2322_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2322_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k2_2322_inst_ack_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2326_inst_req_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2326_inst_ack_0 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2326_inst_req_1 : boolean;
  signal RPIPE_xxconvolvexxconv_k3_2326_inst_ack_1 : boolean;
  signal W_read_k_2284_delayed_1_0_2328_inst_req_0 : boolean;
  signal W_read_k_2284_delayed_1_0_2328_inst_ack_0 : boolean;
  signal W_read_k_2284_delayed_1_0_2328_inst_req_1 : boolean;
  signal W_read_k_2284_delayed_1_0_2328_inst_ack_1 : boolean;
  signal W_read_k_2290_delayed_1_0_2337_inst_req_0 : boolean;
  signal W_read_k_2290_delayed_1_0_2337_inst_ack_0 : boolean;
  signal W_read_k_2290_delayed_1_0_2337_inst_req_1 : boolean;
  signal W_read_k_2290_delayed_1_0_2337_inst_ack_1 : boolean;
  signal W_read_k_2296_delayed_1_0_2346_inst_req_0 : boolean;
  signal W_read_k_2296_delayed_1_0_2346_inst_ack_0 : boolean;
  signal W_read_k_2296_delayed_1_0_2346_inst_req_1 : boolean;
  signal W_read_k_2296_delayed_1_0_2346_inst_ack_1 : boolean;
  signal slice_2357_inst_req_0 : boolean;
  signal slice_2357_inst_ack_0 : boolean;
  signal slice_2357_inst_req_1 : boolean;
  signal slice_2357_inst_ack_1 : boolean;
  signal slice_2361_inst_req_0 : boolean;
  signal slice_2361_inst_ack_0 : boolean;
  signal slice_2361_inst_req_1 : boolean;
  signal slice_2361_inst_ack_1 : boolean;
  signal slice_2365_inst_req_0 : boolean;
  signal slice_2365_inst_ack_0 : boolean;
  signal slice_2365_inst_req_1 : boolean;
  signal slice_2365_inst_ack_1 : boolean;
  signal slice_2369_inst_req_0 : boolean;
  signal slice_2369_inst_ack_0 : boolean;
  signal slice_2369_inst_req_1 : boolean;
  signal slice_2369_inst_ack_1 : boolean;
  signal slice_2373_inst_req_0 : boolean;
  signal slice_2373_inst_ack_0 : boolean;
  signal slice_2373_inst_req_1 : boolean;
  signal slice_2373_inst_ack_1 : boolean;
  signal slice_2377_inst_req_0 : boolean;
  signal slice_2377_inst_ack_0 : boolean;
  signal slice_2377_inst_req_1 : boolean;
  signal slice_2377_inst_ack_1 : boolean;
  signal slice_2381_inst_req_0 : boolean;
  signal slice_2381_inst_ack_0 : boolean;
  signal slice_2381_inst_req_1 : boolean;
  signal slice_2381_inst_ack_1 : boolean;
  signal slice_2385_inst_req_0 : boolean;
  signal slice_2385_inst_ack_0 : boolean;
  signal slice_2385_inst_req_1 : boolean;
  signal slice_2385_inst_ack_1 : boolean;
  signal slice_2389_inst_req_0 : boolean;
  signal slice_2389_inst_ack_0 : boolean;
  signal slice_2389_inst_req_1 : boolean;
  signal slice_2389_inst_ack_1 : boolean;
  signal slice_2393_inst_req_0 : boolean;
  signal slice_2393_inst_ack_0 : boolean;
  signal slice_2393_inst_req_1 : boolean;
  signal slice_2393_inst_ack_1 : boolean;
  signal W_store_kernel_2945_delayed_1_0_3011_inst_req_0 : boolean;
  signal W_store_kernel_2945_delayed_1_0_3011_inst_ack_0 : boolean;
  signal W_store_kernel_2945_delayed_1_0_3011_inst_req_1 : boolean;
  signal W_store_kernel_2945_delayed_1_0_3011_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3015_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3015_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3015_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k2_3015_inst_ack_1 : boolean;
  signal W_store_kernel_2949_delayed_1_0_3018_inst_req_0 : boolean;
  signal W_store_kernel_2949_delayed_1_0_3018_inst_ack_0 : boolean;
  signal W_store_kernel_2949_delayed_1_0_3018_inst_req_1 : boolean;
  signal W_store_kernel_2949_delayed_1_0_3018_inst_ack_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3022_inst_req_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3022_inst_ack_0 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3022_inst_req_1 : boolean;
  signal WPIPE_xxconvolvexxconv_k3_3022_inst_ack_1 : boolean;
  signal W_num_done_2992_delayed_2_0_3063_inst_req_0 : boolean;
  signal W_num_done_2992_delayed_2_0_3063_inst_ack_0 : boolean;
  signal W_num_done_2992_delayed_2_0_3063_inst_req_1 : boolean;
  signal W_num_done_2992_delayed_2_0_3063_inst_ack_1 : boolean;
  signal W_num_done_2998_delayed_2_0_3072_inst_req_0 : boolean;
  signal W_num_done_2998_delayed_2_0_3072_inst_ack_0 : boolean;
  signal W_num_done_2998_delayed_2_0_3072_inst_req_1 : boolean;
  signal W_num_done_2998_delayed_2_0_3072_inst_ack_1 : boolean;
  signal W_num_done_3003_delayed_2_0_3081_inst_req_0 : boolean;
  signal W_num_done_3003_delayed_2_0_3081_inst_ack_0 : boolean;
  signal W_num_done_3003_delayed_2_0_3081_inst_req_1 : boolean;
  signal W_num_done_3003_delayed_2_0_3081_inst_ack_1 : boolean;
  signal CONCAT_u8_u16_3090_inst_req_0 : boolean;
  signal CONCAT_u8_u16_3090_inst_ack_0 : boolean;
  signal CONCAT_u8_u16_3090_inst_req_1 : boolean;
  signal CONCAT_u8_u16_3090_inst_ack_1 : boolean;
  signal WPIPE_output_pipe_3085_inst_req_0 : boolean;
  signal WPIPE_output_pipe_3085_inst_ack_0 : boolean;
  signal WPIPE_output_pipe_3085_inst_req_1 : boolean;
  signal WPIPE_output_pipe_3085_inst_ack_1 : boolean;
  signal do_while_stmt_1890_branch_ack_0 : boolean;
  signal do_while_stmt_1890_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3095_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3095_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3095_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3095_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convolve_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convolve_CP_4675_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convolve_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4675_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convolve_CP_4675_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convolve_CP_4675_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convolve_CP_4675: Block -- control-path 
    signal convolve_CP_4675_elements: BooleanArray(536 downto 0);
    -- 
  begin -- 
    convolve_CP_4675_elements(0) <= convolve_CP_4675_start;
    convolve_CP_4675_symbol <= convolve_CP_4675_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	536 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1873/$entry
      -- CP-element group 0: 	 branch_block_stmt_1873/branch_block_stmt_1873__entry__
      -- CP-element group 0: 	 branch_block_stmt_1873/merge_stmt_1874__entry__
      -- CP-element group 0: 	 branch_block_stmt_1873/merge_stmt_1874_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1873/merge_stmt_1874__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1873/merge_stmt_1874__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1873/$exit
      -- CP-element group 1: 	 branch_block_stmt_1873/branch_block_stmt_1873__exit__
      -- 
    convolve_CP_4675_elements(1) <= false; 
    -- CP-element group 2:  transition  place  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	533 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	534 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_1873/do_while_stmt_1890__exit__
      -- CP-element group 2: 	 branch_block_stmt_1873/assign_stmt_3097__entry__
      -- CP-element group 2: 	 branch_block_stmt_1873/assign_stmt_3097/$entry
      -- CP-element group 2: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Sample/req
      -- 
    req_6469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(2), ack => WPIPE_input_done_pipe_3095_inst_req_0); -- 
    convolve_CP_4675_elements(2) <= convolve_CP_4675_elements(533);
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	536 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Update/cr
      -- 
    ra_4707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1876_inst_ack_0, ack => convolve_CP_4675_elements(3)); -- 
    cr_4711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(3), ack => RPIPE_num_out_pipe_1876_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Sample/rr
      -- 
    ca_4712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1876_inst_ack_1, ack => convolve_CP_4675_elements(4)); -- 
    rr_4734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(4), ack => RPIPE_num_out_pipe_1881_inst_req_0); -- 
    rr_4716_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4716_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(4), ack => SUB_u16_u16_1878_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Sample/ra
      -- 
    ra_4717_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1878_inst_ack_0, ack => convolve_CP_4675_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	536 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	15 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Update/ca
      -- 
    ca_4722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1878_inst_ack_1, ack => convolve_CP_4675_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_update_start_
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Update/cr
      -- 
    ra_4735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1881_inst_ack_0, ack => convolve_CP_4675_elements(7)); -- 
    cr_4739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(7), ack => RPIPE_num_out_pipe_1881_inst_req_1); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1881_Update/ca
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Sample/rr
      -- 
    ca_4740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_num_out_pipe_1881_inst_ack_1, ack => convolve_CP_4675_elements(8)); -- 
    rr_4744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(8), ack => SUB_u16_u16_1883_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Sample/ra
      -- 
    ra_4745_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1883_inst_ack_0, ack => convolve_CP_4675_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	536 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Update/ca
      -- 
    ca_4750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1883_inst_ack_1, ack => convolve_CP_4675_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	536 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Update/cr
      -- 
    ra_4763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1886_inst_ack_0, ack => convolve_CP_4675_elements(11)); -- 
    cr_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(11), ack => RPIPE_size_pipe_1886_inst_req_1); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Sample/rr
      -- 
    ca_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_size_pipe_1886_inst_ack_1, ack => convolve_CP_4675_elements(12)); -- 
    rr_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(12), ack => SUB_u16_u16_1888_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Sample/ra
      -- 
    ra_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1888_inst_ack_0, ack => convolve_CP_4675_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	536 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Update/ca
      -- 
    ca_4778_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_1888_inst_ack_1, ack => convolve_CP_4675_elements(14)); -- 
    -- CP-element group 15:  join  transition  place  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	6 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889__exit__
      -- CP-element group 15: 	 branch_block_stmt_1873/do_while_stmt_1890__entry__
      -- CP-element group 15: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/$exit
      -- 
    convolve_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(6) & convolve_CP_4675_elements(14) & convolve_CP_4675_elements(10);
      gj_convolve_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	22 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1873/do_while_stmt_1890/$entry
      -- CP-element group 16: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890__entry__
      -- 
    convolve_CP_4675_elements(16) <= convolve_CP_4675_elements(15);
    -- CP-element group 17:  merge  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	533 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890__exit__
      -- 
    -- Element group convolve_CP_4675_elements(17) is bound as output of CP function.
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_back
      -- 
    -- Element group convolve_CP_4675_elements(18) is bound as output of CP function.
    -- CP-element group 19:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	531 
    -- CP-element group 19: 	532 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1873/do_while_stmt_1890/condition_done
      -- CP-element group 19: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_exit/$entry
      -- CP-element group 19: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_taken/$entry
      -- 
    convolve_CP_4675_elements(19) <= convolve_CP_4675_elements(24);
    -- CP-element group 20:  branch  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	530 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_body_done
      -- 
    convolve_CP_4675_elements(20) <= convolve_CP_4675_elements(530);
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	109 
    -- CP-element group 21: 	92 
    -- CP-element group 21: 	73 
    -- CP-element group 21: 	54 
    -- CP-element group 21: 	128 
    -- CP-element group 21: 	35 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/back_edge_to_loop_body
      -- 
    convolve_CP_4675_elements(21) <= convolve_CP_4675_elements(18);
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	111 
    -- CP-element group 22: 	94 
    -- CP-element group 22: 	75 
    -- CP-element group 22: 	130 
    -- CP-element group 22: 	56 
    -- CP-element group 22: 	37 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/first_time_through_loop_body
      -- 
    convolve_CP_4675_elements(22) <= convolve_CP_4675_elements(16);
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	157 
    -- CP-element group 23: 	161 
    -- CP-element group 23: 	105 
    -- CP-element group 23: 	106 
    -- CP-element group 23: 	345 
    -- CP-element group 23: 	349 
    -- CP-element group 23: 	141 
    -- CP-element group 23: 	357 
    -- CP-element group 23: 	361 
    -- CP-element group 23: 	353 
    -- CP-element group 23: 	48 
    -- CP-element group 23: 	49 
    -- CP-element group 23: 	122 
    -- CP-element group 23: 	123 
    -- CP-element group 23: 	145 
    -- CP-element group 23: 	29 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	86 
    -- CP-element group 23: 	87 
    -- CP-element group 23: 	529 
    -- CP-element group 23: 	67 
    -- CP-element group 23: 	68 
    -- CP-element group 23: 	165 
    -- CP-element group 23: 	169 
    -- CP-element group 23: 	485 
    -- CP-element group 23: 	365 
    -- CP-element group 23: 	149 
    -- CP-element group 23: 	153 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/$entry
      -- CP-element group 23: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/loop_body_start
      -- 
    -- Element group convolve_CP_4675_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	108 
    -- CP-element group 24: 	72 
    -- CP-element group 24: 	127 
    -- CP-element group 24: 	28 
    -- CP-element group 24: 	91 
    -- CP-element group 24: 	529 
    -- CP-element group 24: 	488 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/condition_evaluated
      -- 
    condition_evaluated_4793_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_4793_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(24), ack => do_while_stmt_1890_branch_req_0); -- 
    convolve_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(72) & convolve_CP_4675_elements(127) & convolve_CP_4675_elements(28) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(529) & convolve_CP_4675_elements(488);
      gj_convolve_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	105 
    -- CP-element group 25: 	48 
    -- CP-element group 25: 	122 
    -- CP-element group 25: 	29 
    -- CP-element group 25: 	86 
    -- CP-element group 25: 	67 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	69 
    -- CP-element group 25: 	50 
    -- CP-element group 25: 	124 
    -- CP-element group 25: 	31 
    -- CP-element group 25: 	88 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/aggregated_phi_sample_req
      -- 
    convolve_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(105) & convolve_CP_4675_elements(48) & convolve_CP_4675_elements(122) & convolve_CP_4675_elements(29) & convolve_CP_4675_elements(86) & convolve_CP_4675_elements(67) & convolve_CP_4675_elements(28);
      gj_convolve_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	107 
    -- CP-element group 26: 	70 
    -- CP-element group 26: 	51 
    -- CP-element group 26: 	125 
    -- CP-element group 26: 	32 
    -- CP-element group 26: 	89 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	482 
    -- CP-element group 26: 	422 
    -- CP-element group 26: 	462 
    -- CP-element group 26: 	466 
    -- CP-element group 26: 	334 
    -- CP-element group 26: 	318 
    -- CP-element group 26: 	322 
    -- CP-element group 26: 	326 
    -- CP-element group 26: 	330 
    -- CP-element group 26: 	314 
    -- CP-element group 26: 	474 
    -- CP-element group 26: 	478 
    -- CP-element group 26: 	438 
    -- CP-element group 26: 	442 
    -- CP-element group 26: 	450 
    -- CP-element group 26: 	454 
    -- CP-element group 26: 	458 
    -- CP-element group 26: 	338 
    -- CP-element group 26: 	342 
    -- CP-element group 26: 	515 
    -- CP-element group 26: 	282 
    -- CP-element group 26: 	286 
    -- CP-element group 26: 	290 
    -- CP-element group 26: 	306 
    -- CP-element group 26: 	310 
    -- CP-element group 26: 	410 
    -- CP-element group 26: 	250 
    -- CP-element group 26: 	254 
    -- CP-element group 26: 	218 
    -- CP-element group 26: 	222 
    -- CP-element group 26: 	274 
    -- CP-element group 26: 	278 
    -- CP-element group 26: 	446 
    -- CP-element group 26: 	270 
    -- CP-element group 26: 	390 
    -- CP-element group 26: 	382 
    -- CP-element group 26: 	386 
    -- CP-element group 26: 	258 
    -- CP-element group 26: 	238 
    -- CP-element group 26: 	226 
    -- CP-element group 26: 	426 
    -- CP-element group 26: 	430 
    -- CP-element group 26: 	294 
    -- CP-element group 26: 	298 
    -- CP-element group 26: 	302 
    -- CP-element group 26: 	470 
    -- CP-element group 26: 	402 
    -- CP-element group 26: 	406 
    -- CP-element group 26: 	394 
    -- CP-element group 26: 	398 
    -- CP-element group 26: 	511 
    -- CP-element group 26: 	242 
    -- CP-element group 26: 	246 
    -- CP-element group 26: 	230 
    -- CP-element group 26: 	234 
    -- CP-element group 26: 	262 
    -- CP-element group 26: 	266 
    -- CP-element group 26: 	530 
    -- CP-element group 26: 	414 
    -- CP-element group 26: 	418 
    -- CP-element group 26: 	434 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	105 
    -- CP-element group 26: 	48 
    -- CP-element group 26: 	122 
    -- CP-element group 26: 	29 
    -- CP-element group 26: 	86 
    -- CP-element group 26: 	67 
    -- CP-element group 26:  members (7) 
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/aggregated_phi_sample_ack
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_sample_completed_
      -- 
    convolve_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(107) & convolve_CP_4675_elements(70) & convolve_CP_4675_elements(51) & convolve_CP_4675_elements(125) & convolve_CP_4675_elements(32) & convolve_CP_4675_elements(89);
      gj_convolve_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	106 
    -- CP-element group 27: 	49 
    -- CP-element group 27: 	123 
    -- CP-element group 27: 	30 
    -- CP-element group 27: 	87 
    -- CP-element group 27: 	68 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	71 
    -- CP-element group 27: 	52 
    -- CP-element group 27: 	126 
    -- CP-element group 27: 	90 
    -- CP-element group 27: 	33 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/aggregated_phi_update_req
      -- 
    convolve_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(106) & convolve_CP_4675_elements(49) & convolve_CP_4675_elements(123) & convolve_CP_4675_elements(30) & convolve_CP_4675_elements(87) & convolve_CP_4675_elements(68);
      gj_convolve_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(27), clk => clk, reset => reset); --
    end block;
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	108 
    -- CP-element group 28: 	72 
    -- CP-element group 28: 	53 
    -- CP-element group 28: 	127 
    -- CP-element group 28: 	91 
    -- CP-element group 28: 	34 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	24 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/aggregated_phi_update_ack
      -- 
    convolve_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(72) & convolve_CP_4675_elements(53) & convolve_CP_4675_elements(127) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(34);
      gj_convolve_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	23 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	480 
    -- CP-element group 29: 	420 
    -- CP-element group 29: 	460 
    -- CP-element group 29: 	464 
    -- CP-element group 29: 	312 
    -- CP-element group 29: 	472 
    -- CP-element group 29: 	476 
    -- CP-element group 29: 	436 
    -- CP-element group 29: 	440 
    -- CP-element group 29: 	448 
    -- CP-element group 29: 	452 
    -- CP-element group 29: 	456 
    -- CP-element group 29: 	513 
    -- CP-element group 29: 	280 
    -- CP-element group 29: 	284 
    -- CP-element group 29: 	288 
    -- CP-element group 29: 	308 
    -- CP-element group 29: 	408 
    -- CP-element group 29: 	248 
    -- CP-element group 29: 	252 
    -- CP-element group 29: 	220 
    -- CP-element group 29: 	276 
    -- CP-element group 29: 	444 
    -- CP-element group 29: 	268 
    -- CP-element group 29: 	272 
    -- CP-element group 29: 	388 
    -- CP-element group 29: 	392 
    -- CP-element group 29: 	384 
    -- CP-element group 29: 	256 
    -- CP-element group 29: 	260 
    -- CP-element group 29: 	236 
    -- CP-element group 29: 	240 
    -- CP-element group 29: 	224 
    -- CP-element group 29: 	228 
    -- CP-element group 29: 	424 
    -- CP-element group 29: 	428 
    -- CP-element group 29: 	292 
    -- CP-element group 29: 	296 
    -- CP-element group 29: 	300 
    -- CP-element group 29: 	304 
    -- CP-element group 29: 	468 
    -- CP-element group 29: 	400 
    -- CP-element group 29: 	404 
    -- CP-element group 29: 	396 
    -- CP-element group 29: 	244 
    -- CP-element group 29: 	232 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	264 
    -- CP-element group 29: 	412 
    -- CP-element group 29: 	416 
    -- CP-element group 29: 	432 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	25 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_sample_start_
      -- 
    convolve_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 51) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1,40 => 1,41 => 1,42 => 1,43 => 1,44 => 1,45 => 1,46 => 1,47 => 1,48 => 1,49 => 1,50 => 1,51 => 1);
      constant place_markings: IntegerArray(0 to 51)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1,40 => 1,41 => 1,42 => 1,43 => 1,44 => 1,45 => 1,46 => 1,47 => 1,48 => 1,49 => 1,50 => 1,51 => 1);
      constant place_delays: IntegerArray(0 to 51) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0,41 => 0,42 => 0,43 => 0,44 => 0,45 => 0,46 => 0,47 => 1,48 => 0,49 => 0,50 => 0,51 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 52); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(480) & convolve_CP_4675_elements(420) & convolve_CP_4675_elements(460) & convolve_CP_4675_elements(464) & convolve_CP_4675_elements(312) & convolve_CP_4675_elements(472) & convolve_CP_4675_elements(476) & convolve_CP_4675_elements(436) & convolve_CP_4675_elements(440) & convolve_CP_4675_elements(448) & convolve_CP_4675_elements(452) & convolve_CP_4675_elements(456) & convolve_CP_4675_elements(513) & convolve_CP_4675_elements(280) & convolve_CP_4675_elements(284) & convolve_CP_4675_elements(288) & convolve_CP_4675_elements(308) & convolve_CP_4675_elements(408) & convolve_CP_4675_elements(248) & convolve_CP_4675_elements(252) & convolve_CP_4675_elements(220) & convolve_CP_4675_elements(276) & convolve_CP_4675_elements(444) & convolve_CP_4675_elements(268) & convolve_CP_4675_elements(272) & convolve_CP_4675_elements(388) & convolve_CP_4675_elements(392) & convolve_CP_4675_elements(384) & convolve_CP_4675_elements(256) & convolve_CP_4675_elements(260) & convolve_CP_4675_elements(236) & convolve_CP_4675_elements(240) & convolve_CP_4675_elements(224) & convolve_CP_4675_elements(228) & convolve_CP_4675_elements(424) & convolve_CP_4675_elements(428) & convolve_CP_4675_elements(292) & convolve_CP_4675_elements(296) & convolve_CP_4675_elements(300) & convolve_CP_4675_elements(304) & convolve_CP_4675_elements(468) & convolve_CP_4675_elements(400) & convolve_CP_4675_elements(404) & convolve_CP_4675_elements(396) & convolve_CP_4675_elements(244) & convolve_CP_4675_elements(232) & convolve_CP_4675_elements(26) & convolve_CP_4675_elements(264) & convolve_CP_4675_elements(412) & convolve_CP_4675_elements(416) & convolve_CP_4675_elements(432);
      gj_convolve_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 52, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	23 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	479 
    -- CP-element group 30: 	34 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	27 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_update_start_
      -- 
    convolve_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(479) & convolve_CP_4675_elements(34);
      gj_convolve_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	25 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_sample_start__ps
      -- 
    convolve_CP_4675_elements(31) <= convolve_CP_4675_elements(25);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	26 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(32) is bound as output of CP function.
    -- CP-element group 33:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	27 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_update_start__ps
      -- 
    convolve_CP_4675_elements(33) <= convolve_CP_4675_elements(27);
    -- CP-element group 34:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	477 
    -- CP-element group 34: 	28 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	30 
    -- CP-element group 34:  members (2) 
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_update_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(34) is bound as output of CP function.
    -- CP-element group 35:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	21 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_loopback_trigger
      -- 
    convolve_CP_4675_elements(35) <= convolve_CP_4675_elements(21);
    -- CP-element group 36:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (2) 
      -- CP-element group 36: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_loopback_sample_req
      -- CP-element group 36: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_loopback_sample_req_ps
      -- 
    phi_stmt_1892_loopback_sample_req_4808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1892_loopback_sample_req_4808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(36), ack => phi_stmt_1892_req_1); -- 
    -- Element group convolve_CP_4675_elements(36) is bound as output of CP function.
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	22 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_entry_trigger
      -- 
    convolve_CP_4675_elements(37) <= convolve_CP_4675_elements(22);
    -- CP-element group 38:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (2) 
      -- CP-element group 38: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_entry_sample_req
      -- CP-element group 38: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_entry_sample_req_ps
      -- 
    phi_stmt_1892_entry_sample_req_4811_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1892_entry_sample_req_4811_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(38), ack => phi_stmt_1892_req_0); -- 
    -- Element group convolve_CP_4675_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_phi_mux_ack
      -- CP-element group 39: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1892_phi_mux_ack_ps
      -- 
    phi_stmt_1892_phi_mux_ack_4814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1892_ack_0, ack => convolve_CP_4675_elements(39)); -- 
    -- CP-element group 40:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_sample_start__ps
      -- CP-element group 40: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_sample_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_sample_completed_
      -- 
    -- Element group convolve_CP_4675_elements(40) is bound as output of CP function.
    -- CP-element group 41:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_update_start__ps
      -- CP-element group 41: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_update_start_
      -- 
    -- Element group convolve_CP_4675_elements(41) is bound as output of CP function.
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	43 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_update_completed__ps
      -- 
    convolve_CP_4675_elements(42) <= convolve_CP_4675_elements(43);
    -- CP-element group 43:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	42 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1896_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(41), ack => convolve_CP_4675_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (4) 
      -- CP-element group 44: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_sample_start__ps
      -- CP-element group 44: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Sample/req
      -- 
    req_4835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(44), ack => nacc1_3071_1897_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_update_start__ps
      -- CP-element group 45: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_update_start_
      -- CP-element group 45: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Update/req
      -- 
    req_4840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(45), ack => nacc1_3071_1897_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_sample_completed__ps
      -- CP-element group 46: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Sample/ack
      -- 
    ack_4836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_3071_1897_buf_ack_0, ack => convolve_CP_4675_elements(46)); -- 
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_update_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc1_1897_Update/ack
      -- 
    ack_4841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc1_3071_1897_buf_ack_1, ack => convolve_CP_4675_elements(47)); -- 
    -- CP-element group 48:  join  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	23 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	420 
    -- CP-element group 48: 	460 
    -- CP-element group 48: 	464 
    -- CP-element group 48: 	332 
    -- CP-element group 48: 	336 
    -- CP-element group 48: 	320 
    -- CP-element group 48: 	324 
    -- CP-element group 48: 	328 
    -- CP-element group 48: 	312 
    -- CP-element group 48: 	316 
    -- CP-element group 48: 	472 
    -- CP-element group 48: 	476 
    -- CP-element group 48: 	436 
    -- CP-element group 48: 	440 
    -- CP-element group 48: 	448 
    -- CP-element group 48: 	452 
    -- CP-element group 48: 	456 
    -- CP-element group 48: 	344 
    -- CP-element group 48: 	340 
    -- CP-element group 48: 	280 
    -- CP-element group 48: 	284 
    -- CP-element group 48: 	288 
    -- CP-element group 48: 	308 
    -- CP-element group 48: 	408 
    -- CP-element group 48: 	517 
    -- CP-element group 48: 	252 
    -- CP-element group 48: 	276 
    -- CP-element group 48: 	444 
    -- CP-element group 48: 	268 
    -- CP-element group 48: 	272 
    -- CP-element group 48: 	388 
    -- CP-element group 48: 	392 
    -- CP-element group 48: 	384 
    -- CP-element group 48: 	256 
    -- CP-element group 48: 	260 
    -- CP-element group 48: 	424 
    -- CP-element group 48: 	428 
    -- CP-element group 48: 	292 
    -- CP-element group 48: 	296 
    -- CP-element group 48: 	300 
    -- CP-element group 48: 	304 
    -- CP-element group 48: 	468 
    -- CP-element group 48: 	400 
    -- CP-element group 48: 	404 
    -- CP-element group 48: 	396 
    -- CP-element group 48: 	26 
    -- CP-element group 48: 	264 
    -- CP-element group 48: 	484 
    -- CP-element group 48: 	412 
    -- CP-element group 48: 	416 
    -- CP-element group 48: 	432 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	25 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_sample_start_
      -- 
    convolve_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 51) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1,40 => 1,41 => 1,42 => 1,43 => 1,44 => 1,45 => 1,46 => 1,47 => 1,48 => 1,49 => 1,50 => 1,51 => 1);
      constant place_markings: IntegerArray(0 to 51)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1,40 => 1,41 => 1,42 => 1,43 => 1,44 => 1,45 => 1,46 => 1,47 => 1,48 => 1,49 => 1,50 => 1,51 => 1);
      constant place_delays: IntegerArray(0 to 51) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0,41 => 0,42 => 0,43 => 0,44 => 0,45 => 0,46 => 1,47 => 0,48 => 0,49 => 0,50 => 0,51 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 52); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(420) & convolve_CP_4675_elements(460) & convolve_CP_4675_elements(464) & convolve_CP_4675_elements(332) & convolve_CP_4675_elements(336) & convolve_CP_4675_elements(320) & convolve_CP_4675_elements(324) & convolve_CP_4675_elements(328) & convolve_CP_4675_elements(312) & convolve_CP_4675_elements(316) & convolve_CP_4675_elements(472) & convolve_CP_4675_elements(476) & convolve_CP_4675_elements(436) & convolve_CP_4675_elements(440) & convolve_CP_4675_elements(448) & convolve_CP_4675_elements(452) & convolve_CP_4675_elements(456) & convolve_CP_4675_elements(344) & convolve_CP_4675_elements(340) & convolve_CP_4675_elements(280) & convolve_CP_4675_elements(284) & convolve_CP_4675_elements(288) & convolve_CP_4675_elements(308) & convolve_CP_4675_elements(408) & convolve_CP_4675_elements(517) & convolve_CP_4675_elements(252) & convolve_CP_4675_elements(276) & convolve_CP_4675_elements(444) & convolve_CP_4675_elements(268) & convolve_CP_4675_elements(272) & convolve_CP_4675_elements(388) & convolve_CP_4675_elements(392) & convolve_CP_4675_elements(384) & convolve_CP_4675_elements(256) & convolve_CP_4675_elements(260) & convolve_CP_4675_elements(424) & convolve_CP_4675_elements(428) & convolve_CP_4675_elements(292) & convolve_CP_4675_elements(296) & convolve_CP_4675_elements(300) & convolve_CP_4675_elements(304) & convolve_CP_4675_elements(468) & convolve_CP_4675_elements(400) & convolve_CP_4675_elements(404) & convolve_CP_4675_elements(396) & convolve_CP_4675_elements(26) & convolve_CP_4675_elements(264) & convolve_CP_4675_elements(484) & convolve_CP_4675_elements(412) & convolve_CP_4675_elements(416) & convolve_CP_4675_elements(432);
      gj_convolve_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 52, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	23 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	483 
    -- CP-element group 49: 	53 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	27 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_update_start_
      -- 
    convolve_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(483) & convolve_CP_4675_elements(53);
      gj_convolve_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	25 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_sample_start__ps
      -- 
    convolve_CP_4675_elements(50) <= convolve_CP_4675_elements(25);
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	26 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	27 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_update_start__ps
      -- 
    convolve_CP_4675_elements(52) <= convolve_CP_4675_elements(27);
    -- CP-element group 53:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	481 
    -- CP-element group 53: 	28 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	49 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_update_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(53) is bound as output of CP function.
    -- CP-element group 54:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	21 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_loopback_trigger
      -- 
    convolve_CP_4675_elements(54) <= convolve_CP_4675_elements(21);
    -- CP-element group 55:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_loopback_sample_req
      -- CP-element group 55: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_loopback_sample_req_ps
      -- 
    phi_stmt_1898_loopback_sample_req_4852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1898_loopback_sample_req_4852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(55), ack => phi_stmt_1898_req_1); -- 
    -- Element group convolve_CP_4675_elements(55) is bound as output of CP function.
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	22 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_entry_trigger
      -- 
    convolve_CP_4675_elements(56) <= convolve_CP_4675_elements(22);
    -- CP-element group 57:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_entry_sample_req
      -- CP-element group 57: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_entry_sample_req_ps
      -- 
    phi_stmt_1898_entry_sample_req_4855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1898_entry_sample_req_4855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(57), ack => phi_stmt_1898_req_0); -- 
    -- Element group convolve_CP_4675_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_phi_mux_ack
      -- CP-element group 58: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1898_phi_mux_ack_ps
      -- 
    phi_stmt_1898_phi_mux_ack_4858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1898_ack_0, ack => convolve_CP_4675_elements(58)); -- 
    -- CP-element group 59:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_sample_completed__ps
      -- CP-element group 59: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_sample_start_
      -- 
    -- Element group convolve_CP_4675_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_update_start__ps
      -- 
    -- Element group convolve_CP_4675_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_update_completed__ps
      -- 
    convolve_CP_4675_elements(61) <= convolve_CP_4675_elements(62);
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	61 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1901_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(60), ack => convolve_CP_4675_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (4) 
      -- CP-element group 63: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_sample_start__ps
      -- CP-element group 63: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Sample/req
      -- CP-element group 63: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_sample_start_
      -- 
    req_4879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(63), ack => nacc2_3080_1902_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_update_start__ps
      -- CP-element group 64: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Update/req
      -- CP-element group 64: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_update_start_
      -- 
    req_4884_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4884_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(64), ack => nacc2_3080_1902_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_sample_completed__ps
      -- CP-element group 65: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Sample/ack
      -- CP-element group 65: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_sample_completed_
      -- 
    ack_4880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3080_1902_buf_ack_0, ack => convolve_CP_4675_elements(65)); -- 
    -- CP-element group 66:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_update_completed__ps
      -- CP-element group 66: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_nacc2_1902_Update/ack
      -- 
    ack_4885_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nacc2_3080_1902_buf_ack_1, ack => convolve_CP_4675_elements(66)); -- 
    -- CP-element group 67:  join  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	23 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	26 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	25 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_sample_start_
      -- 
    convolve_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(26);
      gj_convolve_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  join  transition  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	23 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	346 
    -- CP-element group 68: 	72 
    -- CP-element group 68: 	358 
    -- CP-element group 68: 	362 
    -- CP-element group 68: 	350 
    -- CP-element group 68: 	354 
    -- CP-element group 68: 	371 
    -- CP-element group 68: 	498 
    -- CP-element group 68: 	505 
    -- CP-element group 68: 	491 
    -- CP-element group 68: 	366 
    -- CP-element group 68: 	375 
    -- CP-element group 68: 	379 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	27 
    -- CP-element group 68:  members (1) 
      -- CP-element group 68: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_update_start_
      -- 
    convolve_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 13) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_markings: IntegerArray(0 to 13)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1);
      constant place_delays: IntegerArray(0 to 13) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 14); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(346) & convolve_CP_4675_elements(72) & convolve_CP_4675_elements(358) & convolve_CP_4675_elements(362) & convolve_CP_4675_elements(350) & convolve_CP_4675_elements(354) & convolve_CP_4675_elements(371) & convolve_CP_4675_elements(498) & convolve_CP_4675_elements(505) & convolve_CP_4675_elements(491) & convolve_CP_4675_elements(366) & convolve_CP_4675_elements(375) & convolve_CP_4675_elements(379);
      gj_convolve_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 14, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	25 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (1) 
      -- CP-element group 69: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_sample_start__ps
      -- 
    convolve_CP_4675_elements(69) <= convolve_CP_4675_elements(25);
    -- CP-element group 70:  join  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	26 
    -- CP-element group 70:  members (1) 
      -- CP-element group 70: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(70) is bound as output of CP function.
    -- CP-element group 71:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	27 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_update_start__ps
      -- 
    convolve_CP_4675_elements(71) <= convolve_CP_4675_elements(27);
    -- CP-element group 72:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	24 
    -- CP-element group 72: 	346 
    -- CP-element group 72: 	358 
    -- CP-element group 72: 	362 
    -- CP-element group 72: 	350 
    -- CP-element group 72: 	354 
    -- CP-element group 72: 	369 
    -- CP-element group 72: 	373 
    -- CP-element group 72: 	496 
    -- CP-element group 72: 	28 
    -- CP-element group 72: 	503 
    -- CP-element group 72: 	489 
    -- CP-element group 72: 	366 
    -- CP-element group 72: 	377 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	68 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_update_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(72) is bound as output of CP function.
    -- CP-element group 73:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	21 
    -- CP-element group 73: successors 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_loopback_trigger
      -- 
    convolve_CP_4675_elements(73) <= convolve_CP_4675_elements(21);
    -- CP-element group 74:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_loopback_sample_req
      -- CP-element group 74: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_loopback_sample_req_ps
      -- 
    phi_stmt_1903_loopback_sample_req_4896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1903_loopback_sample_req_4896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(74), ack => phi_stmt_1903_req_1); -- 
    -- Element group convolve_CP_4675_elements(74) is bound as output of CP function.
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	22 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_entry_trigger
      -- 
    convolve_CP_4675_elements(75) <= convolve_CP_4675_elements(22);
    -- CP-element group 76:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_entry_sample_req
      -- CP-element group 76: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_entry_sample_req_ps
      -- 
    phi_stmt_1903_entry_sample_req_4899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1903_entry_sample_req_4899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(76), ack => phi_stmt_1903_req_0); -- 
    -- Element group convolve_CP_4675_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_phi_mux_ack_ps
      -- CP-element group 77: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1903_phi_mux_ack
      -- 
    phi_stmt_1903_phi_mux_ack_4902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1903_ack_0, ack => convolve_CP_4675_elements(77)); -- 
    -- CP-element group 78:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (4) 
      -- CP-element group 78: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_sample_start__ps
      -- CP-element group 78: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_sample_completed__ps
      -- CP-element group 78: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_sample_start_
      -- 
    -- Element group convolve_CP_4675_elements(78) is bound as output of CP function.
    -- CP-element group 79:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_update_start__ps
      -- CP-element group 79: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_update_start_
      -- 
    -- Element group convolve_CP_4675_elements(79) is bound as output of CP function.
    -- CP-element group 80:  join  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	81 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_update_completed__ps
      -- 
    convolve_CP_4675_elements(80) <= convolve_CP_4675_elements(81);
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	80 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1906_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(79), ack => convolve_CP_4675_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (4) 
      -- CP-element group 82: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_sample_start__ps
      -- CP-element group 82: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Sample/req
      -- 
    req_4923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(82), ack => n_row_3062_1907_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_update_start__ps
      -- CP-element group 83: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_update_start_
      -- CP-element group 83: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Update/req
      -- 
    req_4928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(83), ack => n_row_3062_1907_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_sample_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Sample/ack
      -- 
    ack_4924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3062_1907_buf_ack_0, ack => convolve_CP_4675_elements(84)); -- 
    -- CP-element group 85:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (4) 
      -- CP-element group 85: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_update_completed__ps
      -- CP-element group 85: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_row_1907_Update/ack
      -- 
    ack_4929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3062_1907_buf_ack_1, ack => convolve_CP_4675_elements(85)); -- 
    -- CP-element group 86:  join  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	23 
    -- CP-element group 86: marked-predecessors 
    -- CP-element group 86: 	26 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	25 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_sample_start_
      -- 
    convolve_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(26);
      gj_convolve_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	23 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	154 
    -- CP-element group 87: 	158 
    -- CP-element group 87: 	162 
    -- CP-element group 87: 	175 
    -- CP-element group 87: 	346 
    -- CP-element group 87: 	191 
    -- CP-element group 87: 	198 
    -- CP-element group 87: 	142 
    -- CP-element group 87: 	358 
    -- CP-element group 87: 	362 
    -- CP-element group 87: 	350 
    -- CP-element group 87: 	354 
    -- CP-element group 87: 	371 
    -- CP-element group 87: 	205 
    -- CP-element group 87: 	212 
    -- CP-element group 87: 	498 
    -- CP-element group 87: 	146 
    -- CP-element group 87: 	183 
    -- CP-element group 87: 	187 
    -- CP-element group 87: 	91 
    -- CP-element group 87: 	179 
    -- CP-element group 87: 	505 
    -- CP-element group 87: 	491 
    -- CP-element group 87: 	166 
    -- CP-element group 87: 	170 
    -- CP-element group 87: 	366 
    -- CP-element group 87: 	150 
    -- CP-element group 87: 	375 
    -- CP-element group 87: 	379 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	27 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_update_start_
      -- 
    convolve_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 29) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_markings: IntegerArray(0 to 29)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1);
      constant place_delays: IntegerArray(0 to 29) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0);
      constant joinName: string(1 to 28) := "convolve_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 30); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(154) & convolve_CP_4675_elements(158) & convolve_CP_4675_elements(162) & convolve_CP_4675_elements(175) & convolve_CP_4675_elements(346) & convolve_CP_4675_elements(191) & convolve_CP_4675_elements(198) & convolve_CP_4675_elements(142) & convolve_CP_4675_elements(358) & convolve_CP_4675_elements(362) & convolve_CP_4675_elements(350) & convolve_CP_4675_elements(354) & convolve_CP_4675_elements(371) & convolve_CP_4675_elements(205) & convolve_CP_4675_elements(212) & convolve_CP_4675_elements(498) & convolve_CP_4675_elements(146) & convolve_CP_4675_elements(183) & convolve_CP_4675_elements(187) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(179) & convolve_CP_4675_elements(505) & convolve_CP_4675_elements(491) & convolve_CP_4675_elements(166) & convolve_CP_4675_elements(170) & convolve_CP_4675_elements(366) & convolve_CP_4675_elements(150) & convolve_CP_4675_elements(375) & convolve_CP_4675_elements(379);
      gj_convolve_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 30, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	25 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_sample_start__ps
      -- 
    convolve_CP_4675_elements(88) <= convolve_CP_4675_elements(25);
    -- CP-element group 89:  join  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	26 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(89) is bound as output of CP function.
    -- CP-element group 90:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	27 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_update_start__ps
      -- 
    convolve_CP_4675_elements(90) <= convolve_CP_4675_elements(27);
    -- CP-element group 91:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	154 
    -- CP-element group 91: 	158 
    -- CP-element group 91: 	162 
    -- CP-element group 91: 	24 
    -- CP-element group 91: 	173 
    -- CP-element group 91: 	346 
    -- CP-element group 91: 	189 
    -- CP-element group 91: 	196 
    -- CP-element group 91: 	142 
    -- CP-element group 91: 	358 
    -- CP-element group 91: 	362 
    -- CP-element group 91: 	350 
    -- CP-element group 91: 	354 
    -- CP-element group 91: 	369 
    -- CP-element group 91: 	373 
    -- CP-element group 91: 	203 
    -- CP-element group 91: 	496 
    -- CP-element group 91: 	146 
    -- CP-element group 91: 	185 
    -- CP-element group 91: 	28 
    -- CP-element group 91: 	177 
    -- CP-element group 91: 	181 
    -- CP-element group 91: 	503 
    -- CP-element group 91: 	166 
    -- CP-element group 91: 	170 
    -- CP-element group 91: 	489 
    -- CP-element group 91: 	366 
    -- CP-element group 91: 	150 
    -- CP-element group 91: 	377 
    -- CP-element group 91: 	210 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	87 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_update_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(91) is bound as output of CP function.
    -- CP-element group 92:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	21 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_loopback_trigger
      -- 
    convolve_CP_4675_elements(92) <= convolve_CP_4675_elements(21);
    -- CP-element group 93:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_loopback_sample_req
      -- CP-element group 93: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_loopback_sample_req_ps
      -- 
    phi_stmt_1908_loopback_sample_req_4940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1908_loopback_sample_req_4940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(93), ack => phi_stmt_1908_req_1); -- 
    -- Element group convolve_CP_4675_elements(93) is bound as output of CP function.
    -- CP-element group 94:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	22 
    -- CP-element group 94: successors 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_entry_trigger
      -- 
    convolve_CP_4675_elements(94) <= convolve_CP_4675_elements(22);
    -- CP-element group 95:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_entry_sample_req
      -- CP-element group 95: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_entry_sample_req_ps
      -- 
    phi_stmt_1908_entry_sample_req_4943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1908_entry_sample_req_4943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(95), ack => phi_stmt_1908_req_0); -- 
    -- Element group convolve_CP_4675_elements(95) is bound as output of CP function.
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_phi_mux_ack
      -- CP-element group 96: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1908_phi_mux_ack_ps
      -- 
    phi_stmt_1908_phi_mux_ack_4946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1908_ack_0, ack => convolve_CP_4675_elements(96)); -- 
    -- CP-element group 97:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (4) 
      -- CP-element group 97: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_sample_completed__ps
      -- CP-element group 97: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_sample_start_
      -- CP-element group 97: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_sample_start__ps
      -- 
    -- Element group convolve_CP_4675_elements(97) is bound as output of CP function.
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_update_start__ps
      -- CP-element group 98: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_update_start_
      -- 
    -- Element group convolve_CP_4675_elements(98) is bound as output of CP function.
    -- CP-element group 99:  join  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	100 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_update_completed__ps
      -- 
    convolve_CP_4675_elements(99) <= convolve_CP_4675_elements(100);
    -- CP-element group 100:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	99 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1911_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(100) is a control-delay.
    cp_element_100_delay: control_delay_element  generic map(name => " 100_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(98), ack => convolve_CP_4675_elements(100), clk => clk, reset =>reset);
    -- CP-element group 101:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	103 
    -- CP-element group 101:  members (4) 
      -- CP-element group 101: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_sample_start_
      -- CP-element group 101: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_sample_start__ps
      -- CP-element group 101: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Sample/$entry
      -- CP-element group 101: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Sample/req
      -- 
    req_4967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(101), ack => n_col_3054_1912_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(101) is bound as output of CP function.
    -- CP-element group 102:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (4) 
      -- CP-element group 102: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_update_start_
      -- CP-element group 102: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Update/$entry
      -- CP-element group 102: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Update/req
      -- CP-element group 102: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_update_start__ps
      -- 
    req_4972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(102), ack => n_col_3054_1912_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(102) is bound as output of CP function.
    -- CP-element group 103:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	101 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (4) 
      -- CP-element group 103: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Sample/ack
      -- CP-element group 103: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_sample_completed_
      -- CP-element group 103: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Sample/$exit
      -- CP-element group 103: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_sample_completed__ps
      -- 
    ack_4968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3054_1912_buf_ack_0, ack => convolve_CP_4675_elements(103)); -- 
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (4) 
      -- CP-element group 104: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_update_completed__ps
      -- CP-element group 104: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_update_completed_
      -- CP-element group 104: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Update/$exit
      -- CP-element group 104: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_col_1912_Update/ack
      -- 
    ack_4973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3054_1912_buf_ack_1, ack => convolve_CP_4675_elements(104)); -- 
    -- CP-element group 105:  join  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	23 
    -- CP-element group 105: marked-predecessors 
    -- CP-element group 105: 	26 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	25 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_sample_start_
      -- 
    convolve_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(26);
      gj_convolve_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  join  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	23 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	154 
    -- CP-element group 106: 	158 
    -- CP-element group 106: 	162 
    -- CP-element group 106: 	108 
    -- CP-element group 106: 	175 
    -- CP-element group 106: 	512 
    -- CP-element group 106: 	516 
    -- CP-element group 106: 	191 
    -- CP-element group 106: 	520 
    -- CP-element group 106: 	198 
    -- CP-element group 106: 	142 
    -- CP-element group 106: 	205 
    -- CP-element group 106: 	212 
    -- CP-element group 106: 	146 
    -- CP-element group 106: 	183 
    -- CP-element group 106: 	187 
    -- CP-element group 106: 	179 
    -- CP-element group 106: 	166 
    -- CP-element group 106: 	170 
    -- CP-element group 106: 	150 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	27 
    -- CP-element group 106:  members (1) 
      -- CP-element group 106: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_update_start_
      -- 
    convolve_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 20) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_markings: IntegerArray(0 to 20)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1);
      constant place_delays: IntegerArray(0 to 20) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 21); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(154) & convolve_CP_4675_elements(158) & convolve_CP_4675_elements(162) & convolve_CP_4675_elements(108) & convolve_CP_4675_elements(175) & convolve_CP_4675_elements(512) & convolve_CP_4675_elements(516) & convolve_CP_4675_elements(191) & convolve_CP_4675_elements(520) & convolve_CP_4675_elements(198) & convolve_CP_4675_elements(142) & convolve_CP_4675_elements(205) & convolve_CP_4675_elements(212) & convolve_CP_4675_elements(146) & convolve_CP_4675_elements(183) & convolve_CP_4675_elements(187) & convolve_CP_4675_elements(179) & convolve_CP_4675_elements(166) & convolve_CP_4675_elements(170) & convolve_CP_4675_elements(150);
      gj_convolve_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 21, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	26 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(107) is bound as output of CP function.
    -- CP-element group 108:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	154 
    -- CP-element group 108: 	158 
    -- CP-element group 108: 	162 
    -- CP-element group 108: 	24 
    -- CP-element group 108: 	173 
    -- CP-element group 108: 	514 
    -- CP-element group 108: 	189 
    -- CP-element group 108: 	518 
    -- CP-element group 108: 	196 
    -- CP-element group 108: 	142 
    -- CP-element group 108: 	203 
    -- CP-element group 108: 	510 
    -- CP-element group 108: 	146 
    -- CP-element group 108: 	185 
    -- CP-element group 108: 	28 
    -- CP-element group 108: 	177 
    -- CP-element group 108: 	181 
    -- CP-element group 108: 	166 
    -- CP-element group 108: 	170 
    -- CP-element group 108: 	150 
    -- CP-element group 108: 	210 
    -- CP-element group 108: marked-successors 
    -- CP-element group 108: 	106 
    -- CP-element group 108:  members (2) 
      -- CP-element group 108: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_update_completed_
      -- CP-element group 108: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_update_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(108) is bound as output of CP function.
    -- CP-element group 109:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	21 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (1) 
      -- CP-element group 109: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_loopback_trigger
      -- 
    convolve_CP_4675_elements(109) <= convolve_CP_4675_elements(21);
    -- CP-element group 110:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_loopback_sample_req_ps
      -- CP-element group 110: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_loopback_sample_req
      -- 
    phi_stmt_1913_loopback_sample_req_4984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1913_loopback_sample_req_4984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(110), ack => phi_stmt_1913_req_1); -- 
    -- Element group convolve_CP_4675_elements(110) is bound as output of CP function.
    -- CP-element group 111:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	22 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_entry_trigger
      -- 
    convolve_CP_4675_elements(111) <= convolve_CP_4675_elements(22);
    -- CP-element group 112:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (2) 
      -- CP-element group 112: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_entry_sample_req
      -- CP-element group 112: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_entry_sample_req_ps
      -- 
    phi_stmt_1913_entry_sample_req_4987_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1913_entry_sample_req_4987_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(112), ack => phi_stmt_1913_req_0); -- 
    -- Element group convolve_CP_4675_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_phi_mux_ack_ps
      -- CP-element group 113: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1913_phi_mux_ack
      -- 
    phi_stmt_1913_phi_mux_ack_4990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1913_ack_0, ack => convolve_CP_4675_elements(113)); -- 
    -- CP-element group 114:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_sample_start__ps
      -- CP-element group 114: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_sample_completed__ps
      -- CP-element group 114: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_sample_completed_
      -- 
    -- Element group convolve_CP_4675_elements(114) is bound as output of CP function.
    -- CP-element group 115:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (2) 
      -- CP-element group 115: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_update_start__ps
      -- CP-element group 115: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_update_start_
      -- 
    -- Element group convolve_CP_4675_elements(115) is bound as output of CP function.
    -- CP-element group 116:  join  transition  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	117 
    -- CP-element group 116: successors 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_update_completed__ps
      -- 
    convolve_CP_4675_elements(116) <= convolve_CP_4675_elements(117);
    -- CP-element group 117:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	116 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1917_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(115), ack => convolve_CP_4675_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (4) 
      -- CP-element group 118: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_sample_start_
      -- CP-element group 118: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_sample_start__ps
      -- CP-element group 118: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Sample/$entry
      -- CP-element group 118: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Sample/req
      -- 
    req_5011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(118), ack => n_num_3043_1918_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(118) is bound as output of CP function.
    -- CP-element group 119:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (4) 
      -- CP-element group 119: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_update_start__ps
      -- CP-element group 119: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Update/$entry
      -- CP-element group 119: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Update/req
      -- CP-element group 119: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_update_start_
      -- 
    req_5016_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5016_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(119), ack => n_num_3043_1918_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(119) is bound as output of CP function.
    -- CP-element group 120:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120:  members (4) 
      -- CP-element group 120: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_sample_completed__ps
      -- CP-element group 120: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Sample/ack
      -- CP-element group 120: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_sample_completed_
      -- CP-element group 120: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Sample/$exit
      -- 
    ack_5012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_3043_1918_buf_ack_0, ack => convolve_CP_4675_elements(120)); -- 
    -- CP-element group 121:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121:  members (4) 
      -- CP-element group 121: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_update_completed__ps
      -- CP-element group 121: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Update/$exit
      -- CP-element group 121: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_Update/ack
      -- CP-element group 121: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_num_1918_update_completed_
      -- 
    ack_5017_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_num_3043_1918_buf_ack_1, ack => convolve_CP_4675_elements(121)); -- 
    -- CP-element group 122:  join  transition  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	23 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	26 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	25 
    -- CP-element group 122:  members (1) 
      -- CP-element group 122: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_sample_start_
      -- 
    convolve_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(26);
      gj_convolve_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  join  transition  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	23 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	512 
    -- CP-element group 123: 	516 
    -- CP-element group 123: 	520 
    -- CP-element group 123: 	127 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	27 
    -- CP-element group 123:  members (1) 
      -- CP-element group 123: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_update_start_
      -- 
    convolve_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(512) & convolve_CP_4675_elements(516) & convolve_CP_4675_elements(520) & convolve_CP_4675_elements(127);
      gj_convolve_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	25 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (1) 
      -- CP-element group 124: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_sample_start__ps
      -- 
    convolve_CP_4675_elements(124) <= convolve_CP_4675_elements(25);
    -- CP-element group 125:  join  transition  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	26 
    -- CP-element group 125:  members (1) 
      -- CP-element group 125: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(125) is bound as output of CP function.
    -- CP-element group 126:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	27 
    -- CP-element group 126: successors 
    -- CP-element group 126:  members (1) 
      -- CP-element group 126: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_update_start__ps
      -- 
    convolve_CP_4675_elements(126) <= convolve_CP_4675_elements(27);
    -- CP-element group 127:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	24 
    -- CP-element group 127: 	514 
    -- CP-element group 127: 	518 
    -- CP-element group 127: 	510 
    -- CP-element group 127: 	28 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	123 
    -- CP-element group 127:  members (2) 
      -- CP-element group 127: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_update_completed__ps
      -- CP-element group 127: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(127) is bound as output of CP function.
    -- CP-element group 128:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	21 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (1) 
      -- CP-element group 128: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_loopback_trigger
      -- 
    convolve_CP_4675_elements(128) <= convolve_CP_4675_elements(21);
    -- CP-element group 129:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: successors 
    -- CP-element group 129:  members (2) 
      -- CP-element group 129: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_loopback_sample_req_ps
      -- CP-element group 129: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_loopback_sample_req
      -- 
    phi_stmt_1919_loopback_sample_req_5028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1919_loopback_sample_req_5028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(129), ack => phi_stmt_1919_req_1); -- 
    -- Element group convolve_CP_4675_elements(129) is bound as output of CP function.
    -- CP-element group 130:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	22 
    -- CP-element group 130: successors 
    -- CP-element group 130:  members (1) 
      -- CP-element group 130: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_entry_trigger
      -- 
    convolve_CP_4675_elements(130) <= convolve_CP_4675_elements(22);
    -- CP-element group 131:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: successors 
    -- CP-element group 131:  members (2) 
      -- CP-element group 131: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_entry_sample_req
      -- CP-element group 131: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_entry_sample_req_ps
      -- 
    phi_stmt_1919_entry_sample_req_5031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1919_entry_sample_req_5031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(131), ack => phi_stmt_1919_req_0); -- 
    -- Element group convolve_CP_4675_elements(131) is bound as output of CP function.
    -- CP-element group 132:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (2) 
      -- CP-element group 132: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_phi_mux_ack
      -- CP-element group 132: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/phi_stmt_1919_phi_mux_ack_ps
      -- 
    phi_stmt_1919_phi_mux_ack_5034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1919_ack_0, ack => convolve_CP_4675_elements(132)); -- 
    -- CP-element group 133:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: successors 
    -- CP-element group 133:  members (4) 
      -- CP-element group 133: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_sample_start_
      -- CP-element group 133: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_sample_start__ps
      -- CP-element group 133: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_sample_completed__ps
      -- 
    -- Element group convolve_CP_4675_elements(133) is bound as output of CP function.
    -- CP-element group 134:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	136 
    -- CP-element group 134:  members (2) 
      -- CP-element group 134: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_update_start__ps
      -- CP-element group 134: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_update_start_
      -- 
    -- Element group convolve_CP_4675_elements(134) is bound as output of CP function.
    -- CP-element group 135:  join  transition  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: successors 
    -- CP-element group 135:  members (1) 
      -- CP-element group 135: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_update_completed__ps
      -- 
    convolve_CP_4675_elements(135) <= convolve_CP_4675_elements(136);
    -- CP-element group 136:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	134 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	135 
    -- CP-element group 136:  members (1) 
      -- CP-element group 136: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/type_cast_1922_update_completed_
      -- 
    -- Element group convolve_CP_4675_elements(136) is a control-delay.
    cp_element_136_delay: control_delay_element  generic map(name => " 136_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(134), ack => convolve_CP_4675_elements(136), clk => clk, reset =>reset);
    -- CP-element group 137:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (4) 
      -- CP-element group 137: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_sample_start__ps
      -- CP-element group 137: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Sample/$entry
      -- CP-element group 137: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Sample/req
      -- CP-element group 137: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_sample_start_
      -- 
    req_5055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(137), ack => n_chl_3032_1923_buf_req_0); -- 
    -- Element group convolve_CP_4675_elements(137) is bound as output of CP function.
    -- CP-element group 138:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	140 
    -- CP-element group 138:  members (4) 
      -- CP-element group 138: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_update_start__ps
      -- CP-element group 138: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_update_start_
      -- CP-element group 138: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Update/req
      -- 
    req_5060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(138), ack => n_chl_3032_1923_buf_req_1); -- 
    -- Element group convolve_CP_4675_elements(138) is bound as output of CP function.
    -- CP-element group 139:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139:  members (4) 
      -- CP-element group 139: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Sample/ack
      -- CP-element group 139: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Sample/$exit
      -- CP-element group 139: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_sample_completed__ps
      -- CP-element group 139: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_sample_completed_
      -- 
    ack_5056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3032_1923_buf_ack_0, ack => convolve_CP_4675_elements(139)); -- 
    -- CP-element group 140:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	138 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (4) 
      -- CP-element group 140: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_update_completed_
      -- CP-element group 140: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_update_completed__ps
      -- CP-element group 140: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Update/$exit
      -- CP-element group 140: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/R_n_chl_1923_Update/ack
      -- 
    ack_5061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3032_1923_buf_ack_1, ack => convolve_CP_4675_elements(140)); -- 
    -- CP-element group 141:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	23 
    -- CP-element group 141: marked-predecessors 
    -- CP-element group 141: 	144 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	143 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_sample_start_
      -- CP-element group 141: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Sample/$entry
      -- CP-element group 141: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Sample/rr
      -- 
    rr_5070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(141), ack => RPIPE_input_pipe1_1936_inst_req_0); -- 
    convolve_cp_element_group_141: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_141"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(144);
      gj_convolve_cp_element_group_141 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(141), clk => clk, reset => reset); --
    end block;
    -- CP-element group 142:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	108 
    -- CP-element group 142: 	143 
    -- CP-element group 142: 	91 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	219 
    -- CP-element group 142: 	194 
    -- CP-element group 142: 	239 
    -- CP-element group 142: 	223 
    -- CP-element group 142: 	227 
    -- CP-element group 142: 	243 
    -- CP-element group 142: 	247 
    -- CP-element group 142: 	231 
    -- CP-element group 142: 	235 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	106 
    -- CP-element group 142: 	87 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_update_start_
      -- CP-element group 142: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Update/cr
      -- 
    cr_5075_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5075_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(142), ack => RPIPE_input_pipe1_1936_inst_req_1); -- 
    convolve_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(143) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(219) & convolve_CP_4675_elements(194) & convolve_CP_4675_elements(239) & convolve_CP_4675_elements(223) & convolve_CP_4675_elements(227) & convolve_CP_4675_elements(243) & convolve_CP_4675_elements(247) & convolve_CP_4675_elements(231) & convolve_CP_4675_elements(235);
      gj_convolve_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  transition  input  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	141 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	142 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_sample_completed_
      -- CP-element group 143: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Sample/$exit
      -- CP-element group 143: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Sample/ra
      -- 
    ra_5071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1936_inst_ack_0, ack => convolve_CP_4675_elements(143)); -- 
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	193 
    -- CP-element group 144: 	217 
    -- CP-element group 144: 	221 
    -- CP-element group 144: 	237 
    -- CP-element group 144: 	241 
    -- CP-element group 144: 	225 
    -- CP-element group 144: 	245 
    -- CP-element group 144: 	229 
    -- CP-element group 144: 	233 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	141 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_update_completed_
      -- CP-element group 144: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Update/$exit
      -- CP-element group 144: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe1_1936_Update/ca
      -- 
    ca_5076_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe1_1936_inst_ack_1, ack => convolve_CP_4675_elements(144)); -- 
    -- CP-element group 145:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	23 
    -- CP-element group 145: marked-predecessors 
    -- CP-element group 145: 	148 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	147 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_sample_start_
      -- CP-element group 145: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Sample/$entry
      -- CP-element group 145: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Sample/rr
      -- 
    rr_5084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(145), ack => RPIPE_input_pipe2_1940_inst_req_0); -- 
    convolve_cp_element_group_145: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_145"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(148);
      gj_convolve_cp_element_group_145 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(145), clk => clk, reset => reset); --
    end block;
    -- CP-element group 146:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	108 
    -- CP-element group 146: 	147 
    -- CP-element group 146: 	91 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	251 
    -- CP-element group 146: 	275 
    -- CP-element group 146: 	279 
    -- CP-element group 146: 	267 
    -- CP-element group 146: 	271 
    -- CP-element group 146: 	255 
    -- CP-element group 146: 	259 
    -- CP-element group 146: 	201 
    -- CP-element group 146: 	263 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146: marked-successors 
    -- CP-element group 146: 	106 
    -- CP-element group 146: 	87 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_update_start_
      -- CP-element group 146: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Update/cr
      -- 
    cr_5089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(146), ack => RPIPE_input_pipe2_1940_inst_req_1); -- 
    convolve_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(147) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(251) & convolve_CP_4675_elements(275) & convolve_CP_4675_elements(279) & convolve_CP_4675_elements(267) & convolve_CP_4675_elements(271) & convolve_CP_4675_elements(255) & convolve_CP_4675_elements(259) & convolve_CP_4675_elements(201) & convolve_CP_4675_elements(263);
      gj_convolve_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  transition  input  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	145 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	146 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_sample_completed_
      -- CP-element group 147: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Sample/$exit
      -- CP-element group 147: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Sample/ra
      -- 
    ra_5085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_1940_inst_ack_0, ack => convolve_CP_4675_elements(147)); -- 
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	249 
    -- CP-element group 148: 	253 
    -- CP-element group 148: 	200 
    -- CP-element group 148: 	277 
    -- CP-element group 148: 	269 
    -- CP-element group 148: 	273 
    -- CP-element group 148: 	257 
    -- CP-element group 148: 	261 
    -- CP-element group 148: 	265 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	145 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_update_completed_
      -- CP-element group 148: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Update/$exit
      -- CP-element group 148: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe2_1940_Update/ca
      -- 
    ca_5090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe2_1940_inst_ack_1, ack => convolve_CP_4675_elements(148)); -- 
    -- CP-element group 149:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	23 
    -- CP-element group 149: marked-predecessors 
    -- CP-element group 149: 	152 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	151 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_sample_start_
      -- CP-element group 149: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Sample/$entry
      -- CP-element group 149: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Sample/rr
      -- 
    rr_5098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(149), ack => RPIPE_input_pipe3_1944_inst_req_0); -- 
    convolve_cp_element_group_149: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_149"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(152);
      gj_convolve_cp_element_group_149 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(149), clk => clk, reset => reset); --
    end block;
    -- CP-element group 150:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	108 
    -- CP-element group 150: 	91 
    -- CP-element group 150: 	151 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	283 
    -- CP-element group 150: 	287 
    -- CP-element group 150: 	291 
    -- CP-element group 150: 	307 
    -- CP-element group 150: 	311 
    -- CP-element group 150: 	295 
    -- CP-element group 150: 	299 
    -- CP-element group 150: 	303 
    -- CP-element group 150: 	208 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150: marked-successors 
    -- CP-element group 150: 	106 
    -- CP-element group 150: 	87 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_update_start_
      -- CP-element group 150: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Update/cr
      -- 
    cr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(150), ack => RPIPE_input_pipe3_1944_inst_req_1); -- 
    convolve_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(151) & convolve_CP_4675_elements(283) & convolve_CP_4675_elements(287) & convolve_CP_4675_elements(291) & convolve_CP_4675_elements(307) & convolve_CP_4675_elements(311) & convolve_CP_4675_elements(295) & convolve_CP_4675_elements(299) & convolve_CP_4675_elements(303) & convolve_CP_4675_elements(208);
      gj_convolve_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  transition  input  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	149 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	150 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_sample_completed_
      -- CP-element group 151: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Sample/$exit
      -- CP-element group 151: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Sample/ra
      -- 
    ra_5099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_1944_inst_ack_0, ack => convolve_CP_4675_elements(151)); -- 
    -- CP-element group 152:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	281 
    -- CP-element group 152: 	285 
    -- CP-element group 152: 	289 
    -- CP-element group 152: 	305 
    -- CP-element group 152: 	309 
    -- CP-element group 152: 	293 
    -- CP-element group 152: 	297 
    -- CP-element group 152: 	301 
    -- CP-element group 152: 	207 
    -- CP-element group 152: marked-successors 
    -- CP-element group 152: 	149 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_update_completed_
      -- CP-element group 152: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Update/$exit
      -- CP-element group 152: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe3_1944_Update/ca
      -- 
    ca_5104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe3_1944_inst_ack_1, ack => convolve_CP_4675_elements(152)); -- 
    -- CP-element group 153:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	23 
    -- CP-element group 153: marked-predecessors 
    -- CP-element group 153: 	156 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	155 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_sample_start_
      -- CP-element group 153: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Sample/$entry
      -- CP-element group 153: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Sample/rr
      -- 
    rr_5112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(153), ack => RPIPE_input_pipe4_1948_inst_req_0); -- 
    convolve_cp_element_group_153: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_153"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(156);
      gj_convolve_cp_element_group_153 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(153), clk => clk, reset => reset); --
    end block;
    -- CP-element group 154:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	155 
    -- CP-element group 154: 	108 
    -- CP-element group 154: 	91 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	331 
    -- CP-element group 154: 	335 
    -- CP-element group 154: 	319 
    -- CP-element group 154: 	323 
    -- CP-element group 154: 	327 
    -- CP-element group 154: 	315 
    -- CP-element group 154: 	343 
    -- CP-element group 154: 	339 
    -- CP-element group 154: 	215 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: marked-successors 
    -- CP-element group 154: 	106 
    -- CP-element group 154: 	87 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_update_start_
      -- CP-element group 154: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Update/cr
      -- 
    cr_5117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(154), ack => RPIPE_input_pipe4_1948_inst_req_1); -- 
    convolve_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(155) & convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(331) & convolve_CP_4675_elements(335) & convolve_CP_4675_elements(319) & convolve_CP_4675_elements(323) & convolve_CP_4675_elements(327) & convolve_CP_4675_elements(315) & convolve_CP_4675_elements(343) & convolve_CP_4675_elements(339) & convolve_CP_4675_elements(215);
      gj_convolve_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  transition  input  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	153 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	154 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_sample_completed_
      -- CP-element group 155: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Sample/$exit
      -- CP-element group 155: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Sample/ra
      -- 
    ra_5113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_1948_inst_ack_0, ack => convolve_CP_4675_elements(155)); -- 
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	333 
    -- CP-element group 156: 	321 
    -- CP-element group 156: 	325 
    -- CP-element group 156: 	329 
    -- CP-element group 156: 	313 
    -- CP-element group 156: 	317 
    -- CP-element group 156: 	337 
    -- CP-element group 156: 	341 
    -- CP-element group 156: 	214 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	153 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_update_completed_
      -- CP-element group 156: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Update/$exit
      -- CP-element group 156: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_input_pipe4_1948_Update/ca
      -- 
    ca_5118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_pipe4_1948_inst_ack_1, ack => convolve_CP_4675_elements(156)); -- 
    -- CP-element group 157:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	23 
    -- CP-element group 157: marked-predecessors 
    -- CP-element group 157: 	160 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	159 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_sample_start_
      -- CP-element group 157: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Sample/$entry
      -- CP-element group 157: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Sample/rr
      -- 
    rr_5126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(157), ack => RPIPE_xxconvolvexxconv_ip1_1952_inst_req_0); -- 
    convolve_cp_element_group_157: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_157"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(160);
      gj_convolve_cp_element_group_157 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(157), clk => clk, reset => reset); --
    end block;
    -- CP-element group 158:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	159 
    -- CP-element group 158: 	108 
    -- CP-element group 158: 	91 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	219 
    -- CP-element group 158: 	194 
    -- CP-element group 158: 	239 
    -- CP-element group 158: 	223 
    -- CP-element group 158: 	227 
    -- CP-element group 158: 	243 
    -- CP-element group 158: 	247 
    -- CP-element group 158: 	231 
    -- CP-element group 158: 	235 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: marked-successors 
    -- CP-element group 158: 	106 
    -- CP-element group 158: 	87 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_update_start_
      -- CP-element group 158: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Update/cr
      -- 
    cr_5131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(158), ack => RPIPE_xxconvolvexxconv_ip1_1952_inst_req_1); -- 
    convolve_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(159) & convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(219) & convolve_CP_4675_elements(194) & convolve_CP_4675_elements(239) & convolve_CP_4675_elements(223) & convolve_CP_4675_elements(227) & convolve_CP_4675_elements(243) & convolve_CP_4675_elements(247) & convolve_CP_4675_elements(231) & convolve_CP_4675_elements(235);
      gj_convolve_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  transition  input  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	157 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	158 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_sample_completed_
      -- CP-element group 159: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Sample/$exit
      -- CP-element group 159: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Sample/ra
      -- 
    ra_5127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_0, ack => convolve_CP_4675_elements(159)); -- 
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	193 
    -- CP-element group 160: 	217 
    -- CP-element group 160: 	221 
    -- CP-element group 160: 	237 
    -- CP-element group 160: 	241 
    -- CP-element group 160: 	225 
    -- CP-element group 160: 	245 
    -- CP-element group 160: 	229 
    -- CP-element group 160: 	233 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	157 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_update_completed_
      -- CP-element group 160: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Update/$exit
      -- CP-element group 160: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip1_1952_Update/ca
      -- 
    ca_5132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_1, ack => convolve_CP_4675_elements(160)); -- 
    -- CP-element group 161:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	23 
    -- CP-element group 161: marked-predecessors 
    -- CP-element group 161: 	164 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	163 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_sample_start_
      -- CP-element group 161: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Sample/$entry
      -- CP-element group 161: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Sample/rr
      -- 
    rr_5140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(161), ack => RPIPE_xxconvolvexxconv_ip2_1956_inst_req_0); -- 
    convolve_cp_element_group_161: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_161"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(164);
      gj_convolve_cp_element_group_161 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(161), clk => clk, reset => reset); --
    end block;
    -- CP-element group 162:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	163 
    -- CP-element group 162: 	108 
    -- CP-element group 162: 	91 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	251 
    -- CP-element group 162: 	275 
    -- CP-element group 162: 	279 
    -- CP-element group 162: 	267 
    -- CP-element group 162: 	271 
    -- CP-element group 162: 	255 
    -- CP-element group 162: 	259 
    -- CP-element group 162: 	201 
    -- CP-element group 162: 	263 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: marked-successors 
    -- CP-element group 162: 	106 
    -- CP-element group 162: 	87 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_update_start_
      -- CP-element group 162: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Update/$entry
      -- CP-element group 162: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Update/cr
      -- 
    cr_5145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(162), ack => RPIPE_xxconvolvexxconv_ip2_1956_inst_req_1); -- 
    convolve_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(163) & convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(251) & convolve_CP_4675_elements(275) & convolve_CP_4675_elements(279) & convolve_CP_4675_elements(267) & convolve_CP_4675_elements(271) & convolve_CP_4675_elements(255) & convolve_CP_4675_elements(259) & convolve_CP_4675_elements(201) & convolve_CP_4675_elements(263);
      gj_convolve_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	161 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	162 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Sample/ra
      -- 
    ra_5141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_0, ack => convolve_CP_4675_elements(163)); -- 
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	249 
    -- CP-element group 164: 	253 
    -- CP-element group 164: 	200 
    -- CP-element group 164: 	277 
    -- CP-element group 164: 	269 
    -- CP-element group 164: 	273 
    -- CP-element group 164: 	257 
    -- CP-element group 164: 	261 
    -- CP-element group 164: 	265 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	161 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip2_1956_Update/ca
      -- 
    ca_5146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_1, ack => convolve_CP_4675_elements(164)); -- 
    -- CP-element group 165:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	23 
    -- CP-element group 165: marked-predecessors 
    -- CP-element group 165: 	168 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_sample_start_
      -- CP-element group 165: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Sample/$entry
      -- CP-element group 165: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Sample/rr
      -- 
    rr_5154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(165), ack => RPIPE_xxconvolvexxconv_ip3_1960_inst_req_0); -- 
    convolve_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(168);
      gj_convolve_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	108 
    -- CP-element group 166: 	91 
    -- CP-element group 166: 	167 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	283 
    -- CP-element group 166: 	287 
    -- CP-element group 166: 	291 
    -- CP-element group 166: 	307 
    -- CP-element group 166: 	311 
    -- CP-element group 166: 	295 
    -- CP-element group 166: 	299 
    -- CP-element group 166: 	303 
    -- CP-element group 166: 	208 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	106 
    -- CP-element group 166: 	87 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_update_start_
      -- CP-element group 166: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Update/$entry
      -- CP-element group 166: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Update/cr
      -- 
    cr_5159_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5159_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(166), ack => RPIPE_xxconvolvexxconv_ip3_1960_inst_req_1); -- 
    convolve_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(167) & convolve_CP_4675_elements(283) & convolve_CP_4675_elements(287) & convolve_CP_4675_elements(291) & convolve_CP_4675_elements(307) & convolve_CP_4675_elements(311) & convolve_CP_4675_elements(295) & convolve_CP_4675_elements(299) & convolve_CP_4675_elements(303) & convolve_CP_4675_elements(208);
      gj_convolve_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  transition  input  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	166 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_sample_completed_
      -- CP-element group 167: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Sample/$exit
      -- CP-element group 167: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Sample/ra
      -- 
    ra_5155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_0, ack => convolve_CP_4675_elements(167)); -- 
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	281 
    -- CP-element group 168: 	285 
    -- CP-element group 168: 	289 
    -- CP-element group 168: 	305 
    -- CP-element group 168: 	309 
    -- CP-element group 168: 	293 
    -- CP-element group 168: 	297 
    -- CP-element group 168: 	301 
    -- CP-element group 168: 	207 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	165 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_update_completed_
      -- CP-element group 168: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Update/$exit
      -- CP-element group 168: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip3_1960_Update/ca
      -- 
    ca_5160_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_1, ack => convolve_CP_4675_elements(168)); -- 
    -- CP-element group 169:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	23 
    -- CP-element group 169: marked-predecessors 
    -- CP-element group 169: 	172 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	171 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_sample_start_
      -- CP-element group 169: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Sample/$entry
      -- CP-element group 169: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Sample/rr
      -- 
    rr_5168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(169), ack => RPIPE_xxconvolvexxconv_ip4_1964_inst_req_0); -- 
    convolve_cp_element_group_169: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_169"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(172);
      gj_convolve_cp_element_group_169 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(169), clk => clk, reset => reset); --
    end block;
    -- CP-element group 170:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	108 
    -- CP-element group 170: 	171 
    -- CP-element group 170: 	91 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	331 
    -- CP-element group 170: 	335 
    -- CP-element group 170: 	319 
    -- CP-element group 170: 	323 
    -- CP-element group 170: 	327 
    -- CP-element group 170: 	315 
    -- CP-element group 170: 	343 
    -- CP-element group 170: 	339 
    -- CP-element group 170: 	215 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: marked-successors 
    -- CP-element group 170: 	106 
    -- CP-element group 170: 	87 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_update_start_
      -- CP-element group 170: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Update/$entry
      -- CP-element group 170: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Update/cr
      -- 
    cr_5173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(170), ack => RPIPE_xxconvolvexxconv_ip4_1964_inst_req_1); -- 
    convolve_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(171) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(331) & convolve_CP_4675_elements(335) & convolve_CP_4675_elements(319) & convolve_CP_4675_elements(323) & convolve_CP_4675_elements(327) & convolve_CP_4675_elements(315) & convolve_CP_4675_elements(343) & convolve_CP_4675_elements(339) & convolve_CP_4675_elements(215);
      gj_convolve_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  transition  input  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	169 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	170 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_sample_completed_
      -- CP-element group 171: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Sample/$exit
      -- CP-element group 171: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Sample/ra
      -- 
    ra_5169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_0, ack => convolve_CP_4675_elements(171)); -- 
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	333 
    -- CP-element group 172: 	321 
    -- CP-element group 172: 	325 
    -- CP-element group 172: 	329 
    -- CP-element group 172: 	313 
    -- CP-element group 172: 	317 
    -- CP-element group 172: 	337 
    -- CP-element group 172: 	341 
    -- CP-element group 172: 	214 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	169 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_update_completed_
      -- CP-element group 172: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Update/$exit
      -- CP-element group 172: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_ip4_1964_Update/ca
      -- 
    ca_5174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_1, ack => convolve_CP_4675_elements(172)); -- 
    -- CP-element group 173:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	108 
    -- CP-element group 173: 	91 
    -- CP-element group 173: marked-predecessors 
    -- CP-element group 173: 	175 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	175 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_sample_start_
      -- CP-element group 173: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Sample/$entry
      -- CP-element group 173: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Sample/req
      -- 
    req_5182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(173), ack => W_read_ip_1946_delayed_1_0_1966_inst_req_0); -- 
    convolve_cp_element_group_173: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_173"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(175);
      gj_convolve_cp_element_group_173 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(173), clk => clk, reset => reset); --
    end block;
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: 	219 
    -- CP-element group 174: 	194 
    -- CP-element group 174: 	239 
    -- CP-element group 174: 	223 
    -- CP-element group 174: 	227 
    -- CP-element group 174: 	243 
    -- CP-element group 174: 	247 
    -- CP-element group 174: 	231 
    -- CP-element group 174: 	235 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_update_start_
      -- CP-element group 174: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Update/req
      -- 
    req_5187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(174), ack => W_read_ip_1946_delayed_1_0_1966_inst_req_1); -- 
    convolve_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(176) & convolve_CP_4675_elements(219) & convolve_CP_4675_elements(194) & convolve_CP_4675_elements(239) & convolve_CP_4675_elements(223) & convolve_CP_4675_elements(227) & convolve_CP_4675_elements(243) & convolve_CP_4675_elements(247) & convolve_CP_4675_elements(231) & convolve_CP_4675_elements(235);
      gj_convolve_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	173 
    -- CP-element group 175: successors 
    -- CP-element group 175: marked-successors 
    -- CP-element group 175: 	106 
    -- CP-element group 175: 	173 
    -- CP-element group 175: 	87 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_sample_completed_
      -- CP-element group 175: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Sample/$exit
      -- CP-element group 175: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Sample/ack
      -- 
    ack_5183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1946_delayed_1_0_1966_inst_ack_0, ack => convolve_CP_4675_elements(175)); -- 
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	193 
    -- CP-element group 176: 	217 
    -- CP-element group 176: 	221 
    -- CP-element group 176: 	237 
    -- CP-element group 176: 	241 
    -- CP-element group 176: 	225 
    -- CP-element group 176: 	245 
    -- CP-element group 176: 	229 
    -- CP-element group 176: 	233 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_update_completed_
      -- CP-element group 176: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Update/$exit
      -- CP-element group 176: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1968_Update/ack
      -- 
    ack_5188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1946_delayed_1_0_1966_inst_ack_1, ack => convolve_CP_4675_elements(176)); -- 
    -- CP-element group 177:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	108 
    -- CP-element group 177: 	91 
    -- CP-element group 177: marked-predecessors 
    -- CP-element group 177: 	179 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	179 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_sample_start_
      -- CP-element group 177: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Sample/$entry
      -- CP-element group 177: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Sample/req
      -- 
    req_5196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(177), ack => W_read_ip_1952_delayed_1_0_1975_inst_req_0); -- 
    convolve_cp_element_group_177: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_177"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(179);
      gj_convolve_cp_element_group_177 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(177), clk => clk, reset => reset); --
    end block;
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	251 
    -- CP-element group 178: 	275 
    -- CP-element group 178: 	279 
    -- CP-element group 178: 	267 
    -- CP-element group 178: 	271 
    -- CP-element group 178: 	255 
    -- CP-element group 178: 	259 
    -- CP-element group 178: 	201 
    -- CP-element group 178: 	263 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_update_start_
      -- CP-element group 178: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Update/req
      -- 
    req_5201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(178), ack => W_read_ip_1952_delayed_1_0_1975_inst_req_1); -- 
    convolve_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(251) & convolve_CP_4675_elements(275) & convolve_CP_4675_elements(279) & convolve_CP_4675_elements(267) & convolve_CP_4675_elements(271) & convolve_CP_4675_elements(255) & convolve_CP_4675_elements(259) & convolve_CP_4675_elements(201) & convolve_CP_4675_elements(263) & convolve_CP_4675_elements(180);
      gj_convolve_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	177 
    -- CP-element group 179: successors 
    -- CP-element group 179: marked-successors 
    -- CP-element group 179: 	106 
    -- CP-element group 179: 	87 
    -- CP-element group 179: 	177 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_sample_completed_
      -- CP-element group 179: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Sample/$exit
      -- CP-element group 179: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Sample/ack
      -- 
    ack_5197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1952_delayed_1_0_1975_inst_ack_0, ack => convolve_CP_4675_elements(179)); -- 
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	249 
    -- CP-element group 180: 	253 
    -- CP-element group 180: 	200 
    -- CP-element group 180: 	277 
    -- CP-element group 180: 	269 
    -- CP-element group 180: 	273 
    -- CP-element group 180: 	257 
    -- CP-element group 180: 	261 
    -- CP-element group 180: 	265 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_update_completed_
      -- CP-element group 180: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Update/$exit
      -- CP-element group 180: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1977_Update/ack
      -- 
    ack_5202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1952_delayed_1_0_1975_inst_ack_1, ack => convolve_CP_4675_elements(180)); -- 
    -- CP-element group 181:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	108 
    -- CP-element group 181: 	91 
    -- CP-element group 181: marked-predecessors 
    -- CP-element group 181: 	183 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	183 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_sample_start_
      -- CP-element group 181: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Sample/$entry
      -- CP-element group 181: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Sample/req
      -- 
    req_5210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(181), ack => W_read_ip_1958_delayed_1_0_1984_inst_req_0); -- 
    convolve_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(183);
      gj_convolve_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	283 
    -- CP-element group 182: 	287 
    -- CP-element group 182: 	291 
    -- CP-element group 182: 	307 
    -- CP-element group 182: 	311 
    -- CP-element group 182: 	295 
    -- CP-element group 182: 	299 
    -- CP-element group 182: 	303 
    -- CP-element group 182: 	184 
    -- CP-element group 182: 	208 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_update_start_
      -- CP-element group 182: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Update/req
      -- 
    req_5215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(182), ack => W_read_ip_1958_delayed_1_0_1984_inst_req_1); -- 
    convolve_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(283) & convolve_CP_4675_elements(287) & convolve_CP_4675_elements(291) & convolve_CP_4675_elements(307) & convolve_CP_4675_elements(311) & convolve_CP_4675_elements(295) & convolve_CP_4675_elements(299) & convolve_CP_4675_elements(303) & convolve_CP_4675_elements(184) & convolve_CP_4675_elements(208);
      gj_convolve_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	181 
    -- CP-element group 183: successors 
    -- CP-element group 183: marked-successors 
    -- CP-element group 183: 	106 
    -- CP-element group 183: 	87 
    -- CP-element group 183: 	181 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_sample_completed_
      -- CP-element group 183: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Sample/$exit
      -- CP-element group 183: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Sample/ack
      -- 
    ack_5211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1958_delayed_1_0_1984_inst_ack_0, ack => convolve_CP_4675_elements(183)); -- 
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	281 
    -- CP-element group 184: 	285 
    -- CP-element group 184: 	289 
    -- CP-element group 184: 	305 
    -- CP-element group 184: 	309 
    -- CP-element group 184: 	293 
    -- CP-element group 184: 	297 
    -- CP-element group 184: 	301 
    -- CP-element group 184: 	207 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_update_completed_
      -- CP-element group 184: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Update/$exit
      -- CP-element group 184: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1986_Update/ack
      -- 
    ack_5216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1958_delayed_1_0_1984_inst_ack_1, ack => convolve_CP_4675_elements(184)); -- 
    -- CP-element group 185:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	108 
    -- CP-element group 185: 	91 
    -- CP-element group 185: marked-predecessors 
    -- CP-element group 185: 	187 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	187 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_sample_start_
      -- CP-element group 185: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Sample/req
      -- 
    req_5224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(185), ack => W_read_ip_1964_delayed_1_0_1993_inst_req_0); -- 
    convolve_cp_element_group_185: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_185"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(187);
      gj_convolve_cp_element_group_185 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(185), clk => clk, reset => reset); --
    end block;
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	331 
    -- CP-element group 186: 	335 
    -- CP-element group 186: 	319 
    -- CP-element group 186: 	323 
    -- CP-element group 186: 	327 
    -- CP-element group 186: 	315 
    -- CP-element group 186: 	343 
    -- CP-element group 186: 	339 
    -- CP-element group 186: 	215 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_update_start_
      -- CP-element group 186: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Update/req
      -- 
    req_5229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(186), ack => W_read_ip_1964_delayed_1_0_1993_inst_req_1); -- 
    convolve_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(331) & convolve_CP_4675_elements(335) & convolve_CP_4675_elements(319) & convolve_CP_4675_elements(323) & convolve_CP_4675_elements(327) & convolve_CP_4675_elements(315) & convolve_CP_4675_elements(343) & convolve_CP_4675_elements(339) & convolve_CP_4675_elements(215) & convolve_CP_4675_elements(188);
      gj_convolve_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	185 
    -- CP-element group 187: successors 
    -- CP-element group 187: marked-successors 
    -- CP-element group 187: 	106 
    -- CP-element group 187: 	185 
    -- CP-element group 187: 	87 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_sample_completed_
      -- CP-element group 187: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Sample/$exit
      -- CP-element group 187: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Sample/ack
      -- 
    ack_5225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1964_delayed_1_0_1993_inst_ack_0, ack => convolve_CP_4675_elements(187)); -- 
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	333 
    -- CP-element group 188: 	321 
    -- CP-element group 188: 	325 
    -- CP-element group 188: 	329 
    -- CP-element group 188: 	313 
    -- CP-element group 188: 	317 
    -- CP-element group 188: 	337 
    -- CP-element group 188: 	341 
    -- CP-element group 188: 	214 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_update_completed_
      -- CP-element group 188: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Update/$exit
      -- CP-element group 188: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_1995_Update/ack
      -- 
    ack_5230_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_ip_1964_delayed_1_0_1993_inst_ack_1, ack => convolve_CP_4675_elements(188)); -- 
    -- CP-element group 189:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	108 
    -- CP-element group 189: 	91 
    -- CP-element group 189: marked-predecessors 
    -- CP-element group 189: 	191 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	191 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_sample_start_
      -- CP-element group 189: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Sample/$entry
      -- CP-element group 189: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Sample/req
      -- 
    req_5238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(189), ack => W_write_input_1978_delayed_1_0_2011_inst_req_0); -- 
    convolve_cp_element_group_189: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_189"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(191);
      gj_convolve_cp_element_group_189 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(189), clk => clk, reset => reset); --
    end block;
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: 	194 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_update_start_
      -- CP-element group 190: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Update/req
      -- 
    req_5243_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5243_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(190), ack => W_write_input_1978_delayed_1_0_2011_inst_req_1); -- 
    convolve_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(192) & convolve_CP_4675_elements(194);
      gj_convolve_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	189 
    -- CP-element group 191: successors 
    -- CP-element group 191: marked-successors 
    -- CP-element group 191: 	106 
    -- CP-element group 191: 	189 
    -- CP-element group 191: 	87 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_sample_completed_
      -- CP-element group 191: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Sample/$exit
      -- CP-element group 191: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Sample/ack
      -- 
    ack_5239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1978_delayed_1_0_2011_inst_ack_0, ack => convolve_CP_4675_elements(191)); -- 
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	193 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_update_completed_
      -- CP-element group 192: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Update/$exit
      -- CP-element group 192: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2013_Update/ack
      -- 
    ack_5244_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1978_delayed_1_0_2011_inst_ack_1, ack => convolve_CP_4675_elements(192)); -- 
    -- CP-element group 193:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	160 
    -- CP-element group 193: 	176 
    -- CP-element group 193: 	192 
    -- CP-element group 193: 	144 
    -- CP-element group 193: marked-predecessors 
    -- CP-element group 193: 	195 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	194 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_sample_start_
      -- CP-element group 193: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Sample/$entry
      -- CP-element group 193: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Sample/req
      -- 
    req_5252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(193), ack => WPIPE_xxconvolvexxconv_ip1_2015_inst_req_0); -- 
    convolve_cp_element_group_193: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_193"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(192) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(195);
      gj_convolve_cp_element_group_193 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(193), clk => clk, reset => reset); --
    end block;
    -- CP-element group 194:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	193 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194: marked-successors 
    -- CP-element group 194: 	158 
    -- CP-element group 194: 	174 
    -- CP-element group 194: 	190 
    -- CP-element group 194: 	142 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_sample_completed_
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_update_start_
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Sample/ack
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Update/req
      -- 
    ack_5253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_0, ack => convolve_CP_4675_elements(194)); -- 
    req_5257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(194), ack => WPIPE_xxconvolvexxconv_ip1_2015_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	530 
    -- CP-element group 195: marked-successors 
    -- CP-element group 195: 	193 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip1_2015_Update/ack
      -- 
    ack_5258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_1, ack => convolve_CP_4675_elements(195)); -- 
    -- CP-element group 196:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	108 
    -- CP-element group 196: 	91 
    -- CP-element group 196: marked-predecessors 
    -- CP-element group 196: 	198 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	198 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_sample_start_
      -- CP-element group 196: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Sample/$entry
      -- CP-element group 196: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Sample/req
      -- 
    req_5266_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5266_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(196), ack => W_write_input_1982_delayed_1_0_2018_inst_req_0); -- 
    convolve_cp_element_group_196: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_196"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(198);
      gj_convolve_cp_element_group_196 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(196), clk => clk, reset => reset); --
    end block;
    -- CP-element group 197:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: marked-predecessors 
    -- CP-element group 197: 	199 
    -- CP-element group 197: 	201 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	199 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_update_start_
      -- CP-element group 197: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Update/$entry
      -- CP-element group 197: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Update/req
      -- 
    req_5271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(197), ack => W_write_input_1982_delayed_1_0_2018_inst_req_1); -- 
    convolve_cp_element_group_197: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_197"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(199) & convolve_CP_4675_elements(201);
      gj_convolve_cp_element_group_197 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(197), clk => clk, reset => reset); --
    end block;
    -- CP-element group 198:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	196 
    -- CP-element group 198: successors 
    -- CP-element group 198: marked-successors 
    -- CP-element group 198: 	106 
    -- CP-element group 198: 	196 
    -- CP-element group 198: 	87 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_sample_completed_
      -- CP-element group 198: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Sample/ack
      -- 
    ack_5267_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1982_delayed_1_0_2018_inst_ack_0, ack => convolve_CP_4675_elements(198)); -- 
    -- CP-element group 199:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	197 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: marked-successors 
    -- CP-element group 199: 	197 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_update_completed_
      -- CP-element group 199: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2020_Update/ack
      -- 
    ack_5272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1982_delayed_1_0_2018_inst_ack_1, ack => convolve_CP_4675_elements(199)); -- 
    -- CP-element group 200:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	164 
    -- CP-element group 200: 	199 
    -- CP-element group 200: 	180 
    -- CP-element group 200: 	148 
    -- CP-element group 200: marked-predecessors 
    -- CP-element group 200: 	202 
    -- CP-element group 200: successors 
    -- CP-element group 200: 	201 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_sample_start_
      -- CP-element group 200: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Sample/$entry
      -- CP-element group 200: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Sample/req
      -- 
    req_5280_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5280_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(200), ack => WPIPE_xxconvolvexxconv_ip2_2022_inst_req_0); -- 
    convolve_cp_element_group_200: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_200"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(199) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(202);
      gj_convolve_cp_element_group_200 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(200), clk => clk, reset => reset); --
    end block;
    -- CP-element group 201:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	200 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	202 
    -- CP-element group 201: marked-successors 
    -- CP-element group 201: 	162 
    -- CP-element group 201: 	197 
    -- CP-element group 201: 	146 
    -- CP-element group 201: 	178 
    -- CP-element group 201:  members (6) 
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_sample_completed_
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_update_start_
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Sample/$exit
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Sample/ack
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Update/$entry
      -- CP-element group 201: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Update/req
      -- 
    ack_5281_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_0, ack => convolve_CP_4675_elements(201)); -- 
    req_5285_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5285_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(201), ack => WPIPE_xxconvolvexxconv_ip2_2022_inst_req_1); -- 
    -- CP-element group 202:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	201 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	530 
    -- CP-element group 202: marked-successors 
    -- CP-element group 202: 	200 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_update_completed_
      -- CP-element group 202: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Update/$exit
      -- CP-element group 202: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip2_2022_Update/ack
      -- 
    ack_5286_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_1, ack => convolve_CP_4675_elements(202)); -- 
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	108 
    -- CP-element group 203: 	91 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	205 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_sample_start_
      -- CP-element group 203: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Sample/req
      -- 
    req_5294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(203), ack => W_write_input_1986_delayed_1_0_2025_inst_req_0); -- 
    convolve_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(205);
      gj_convolve_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: marked-predecessors 
    -- CP-element group 204: 	206 
    -- CP-element group 204: 	208 
    -- CP-element group 204: successors 
    -- CP-element group 204: 	206 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_update_start_
      -- CP-element group 204: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Update/$entry
      -- CP-element group 204: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Update/req
      -- 
    req_5299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(204), ack => W_write_input_1986_delayed_1_0_2025_inst_req_1); -- 
    convolve_cp_element_group_204: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_204"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(206) & convolve_CP_4675_elements(208);
      gj_convolve_cp_element_group_204 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(204), clk => clk, reset => reset); --
    end block;
    -- CP-element group 205:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: marked-successors 
    -- CP-element group 205: 	106 
    -- CP-element group 205: 	203 
    -- CP-element group 205: 	87 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_sample_completed_
      -- CP-element group 205: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Sample/$exit
      -- CP-element group 205: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Sample/ack
      -- 
    ack_5295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1986_delayed_1_0_2025_inst_ack_0, ack => convolve_CP_4675_elements(205)); -- 
    -- CP-element group 206:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	204 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206: marked-successors 
    -- CP-element group 206: 	204 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_update_completed_
      -- CP-element group 206: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Update/$exit
      -- CP-element group 206: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2027_Update/ack
      -- 
    ack_5300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 206_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1986_delayed_1_0_2025_inst_ack_1, ack => convolve_CP_4675_elements(206)); -- 
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	184 
    -- CP-element group 207: 	168 
    -- CP-element group 207: 	152 
    -- CP-element group 207: 	206 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	209 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	208 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_sample_start_
      -- CP-element group 207: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Sample/$entry
      -- CP-element group 207: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Sample/req
      -- 
    req_5308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(207), ack => WPIPE_xxconvolvexxconv_ip3_2029_inst_req_0); -- 
    convolve_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(206) & convolve_CP_4675_elements(209);
      gj_convolve_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	207 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	204 
    -- CP-element group 208: 	182 
    -- CP-element group 208: 	166 
    -- CP-element group 208: 	150 
    -- CP-element group 208:  members (6) 
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_update_start_
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Sample/ack
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Update/$entry
      -- CP-element group 208: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Update/req
      -- 
    ack_5309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_0, ack => convolve_CP_4675_elements(208)); -- 
    req_5313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(208), ack => WPIPE_xxconvolvexxconv_ip3_2029_inst_req_1); -- 
    -- CP-element group 209:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	530 
    -- CP-element group 209: marked-successors 
    -- CP-element group 209: 	207 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip3_2029_Update/ack
      -- 
    ack_5314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_1, ack => convolve_CP_4675_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	108 
    -- CP-element group 210: 	91 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Sample/req
      -- 
    req_5322_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5322_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(210), ack => W_write_input_1990_delayed_1_0_2032_inst_req_0); -- 
    convolve_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(212);
      gj_convolve_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	213 
    -- CP-element group 211: 	215 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_update_start_
      -- CP-element group 211: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Update/req
      -- 
    req_5327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(211), ack => W_write_input_1990_delayed_1_0_2032_inst_req_1); -- 
    convolve_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(213) & convolve_CP_4675_elements(215);
      gj_convolve_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	106 
    -- CP-element group 212: 	87 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Sample/ack
      -- 
    ack_5323_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1990_delayed_1_0_2032_inst_ack_0, ack => convolve_CP_4675_elements(212)); -- 
    -- CP-element group 213:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	214 
    -- CP-element group 213: marked-successors 
    -- CP-element group 213: 	211 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2034_Update/ack
      -- 
    ack_5328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_input_1990_delayed_1_0_2032_inst_ack_1, ack => convolve_CP_4675_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	156 
    -- CP-element group 214: 	172 
    -- CP-element group 214: 	213 
    -- CP-element group 214: 	188 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	215 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Sample/req
      -- 
    req_5336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(214), ack => WPIPE_xxconvolvexxconv_ip4_2036_inst_req_0); -- 
    convolve_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(213) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(216);
      gj_convolve_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	214 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	216 
    -- CP-element group 215: marked-successors 
    -- CP-element group 215: 	154 
    -- CP-element group 215: 	186 
    -- CP-element group 215: 	170 
    -- CP-element group 215: 	211 
    -- CP-element group 215:  members (6) 
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_sample_completed_
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_update_start_
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Sample/$exit
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Sample/ack
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Update/req
      -- 
    ack_5337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_0, ack => convolve_CP_4675_elements(215)); -- 
    req_5341_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5341_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(215), ack => WPIPE_xxconvolvexxconv_ip4_2036_inst_req_1); -- 
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	215 
    -- CP-element group 216: successors 
    -- CP-element group 216: 	530 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_update_completed_
      -- CP-element group 216: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Update/$exit
      -- CP-element group 216: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_ip4_2036_Update/ack
      -- 
    ack_5342_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_1, ack => convolve_CP_4675_elements(216)); -- 
    -- CP-element group 217:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	160 
    -- CP-element group 217: 	176 
    -- CP-element group 217: 	144 
    -- CP-element group 217: marked-predecessors 
    -- CP-element group 217: 	219 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	219 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_sample_start_
      -- CP-element group 217: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Sample/$entry
      -- CP-element group 217: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Sample/rr
      -- 
    rr_5350_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5350_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(217), ack => slice_2041_inst_req_0); -- 
    convolve_cp_element_group_217: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_217"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(219);
      gj_convolve_cp_element_group_217 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(217), clk => clk, reset => reset); --
    end block;
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	26 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: 	524 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_update_start_
      -- CP-element group 218: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Update/$entry
      -- CP-element group 218: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Update/cr
      -- 
    cr_5355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(218), ack => slice_2041_inst_req_1); -- 
    convolve_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(220) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	217 
    -- CP-element group 219: successors 
    -- CP-element group 219: marked-successors 
    -- CP-element group 219: 	158 
    -- CP-element group 219: 	174 
    -- CP-element group 219: 	217 
    -- CP-element group 219: 	142 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_sample_completed_
      -- CP-element group 219: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Sample/$exit
      -- CP-element group 219: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Sample/ra
      -- 
    ra_5351_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2041_inst_ack_0, ack => convolve_CP_4675_elements(219)); -- 
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	522 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: 	29 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_update_completed_
      -- CP-element group 220: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Update/$exit
      -- CP-element group 220: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2041_Update/ca
      -- 
    ca_5356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2041_inst_ack_1, ack => convolve_CP_4675_elements(220)); -- 
    -- CP-element group 221:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	160 
    -- CP-element group 221: 	176 
    -- CP-element group 221: 	144 
    -- CP-element group 221: marked-predecessors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_sample_start_
      -- CP-element group 221: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Sample/$entry
      -- CP-element group 221: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Sample/rr
      -- 
    rr_5364_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5364_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(221), ack => slice_2045_inst_req_0); -- 
    convolve_cp_element_group_221: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_221"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(223);
      gj_convolve_cp_element_group_221 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(221), clk => clk, reset => reset); --
    end block;
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	26 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: 	524 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_update_start_
      -- CP-element group 222: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Update/$entry
      -- CP-element group 222: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Update/cr
      -- 
    cr_5369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(222), ack => slice_2045_inst_req_1); -- 
    convolve_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(224) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	221 
    -- CP-element group 223: successors 
    -- CP-element group 223: marked-successors 
    -- CP-element group 223: 	158 
    -- CP-element group 223: 	174 
    -- CP-element group 223: 	221 
    -- CP-element group 223: 	142 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_sample_completed_
      -- CP-element group 223: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Sample/ra
      -- 
    ra_5365_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2045_inst_ack_0, ack => convolve_CP_4675_elements(223)); -- 
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	522 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: 	29 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_update_completed_
      -- CP-element group 224: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2045_Update/ca
      -- 
    ca_5370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2045_inst_ack_1, ack => convolve_CP_4675_elements(224)); -- 
    -- CP-element group 225:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	160 
    -- CP-element group 225: 	176 
    -- CP-element group 225: 	144 
    -- CP-element group 225: marked-predecessors 
    -- CP-element group 225: 	227 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	227 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_sample_start_
      -- CP-element group 225: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Sample/$entry
      -- CP-element group 225: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Sample/rr
      -- 
    rr_5378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(225), ack => slice_2049_inst_req_0); -- 
    convolve_cp_element_group_225: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_225"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(227);
      gj_convolve_cp_element_group_225 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(225), clk => clk, reset => reset); --
    end block;
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	26 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: 	524 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_update_start_
      -- CP-element group 226: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Update/$entry
      -- CP-element group 226: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Update/cr
      -- 
    cr_5383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(226), ack => slice_2049_inst_req_1); -- 
    convolve_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(228) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	225 
    -- CP-element group 227: successors 
    -- CP-element group 227: marked-successors 
    -- CP-element group 227: 	158 
    -- CP-element group 227: 	174 
    -- CP-element group 227: 	142 
    -- CP-element group 227: 	225 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Sample/ra
      -- 
    ra_5379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2049_inst_ack_0, ack => convolve_CP_4675_elements(227)); -- 
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	522 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	29 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2049_Update/ca
      -- 
    ca_5384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2049_inst_ack_1, ack => convolve_CP_4675_elements(228)); -- 
    -- CP-element group 229:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	160 
    -- CP-element group 229: 	176 
    -- CP-element group 229: 	144 
    -- CP-element group 229: marked-predecessors 
    -- CP-element group 229: 	231 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_sample_start_
      -- CP-element group 229: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Sample/$entry
      -- CP-element group 229: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Sample/rr
      -- 
    rr_5392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(229), ack => slice_2053_inst_req_0); -- 
    convolve_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(231);
      gj_convolve_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	26 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	524 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_update_start_
      -- CP-element group 230: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Update/$entry
      -- CP-element group 230: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Update/cr
      -- 
    cr_5397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(230), ack => slice_2053_inst_req_1); -- 
    convolve_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(232);
      gj_convolve_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: marked-successors 
    -- CP-element group 231: 	158 
    -- CP-element group 231: 	174 
    -- CP-element group 231: 	142 
    -- CP-element group 231: 	229 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_sample_completed_
      -- CP-element group 231: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Sample/$exit
      -- CP-element group 231: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Sample/ra
      -- 
    ra_5393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2053_inst_ack_0, ack => convolve_CP_4675_elements(231)); -- 
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: 	522 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: 	29 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_update_completed_
      -- CP-element group 232: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Update/$exit
      -- CP-element group 232: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2053_Update/ca
      -- 
    ca_5398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2053_inst_ack_1, ack => convolve_CP_4675_elements(232)); -- 
    -- CP-element group 233:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	160 
    -- CP-element group 233: 	176 
    -- CP-element group 233: 	144 
    -- CP-element group 233: marked-predecessors 
    -- CP-element group 233: 	235 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	235 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_sample_start_
      -- CP-element group 233: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Sample/$entry
      -- CP-element group 233: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Sample/rr
      -- 
    rr_5406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(233), ack => slice_2057_inst_req_0); -- 
    convolve_cp_element_group_233: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_233"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(235);
      gj_convolve_cp_element_group_233 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(233), clk => clk, reset => reset); --
    end block;
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	26 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: 	524 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_update_start_
      -- CP-element group 234: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Update/$entry
      -- CP-element group 234: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Update/cr
      -- 
    cr_5411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(234), ack => slice_2057_inst_req_1); -- 
    convolve_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(236) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	233 
    -- CP-element group 235: successors 
    -- CP-element group 235: marked-successors 
    -- CP-element group 235: 	158 
    -- CP-element group 235: 	174 
    -- CP-element group 235: 	142 
    -- CP-element group 235: 	233 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_sample_completed_
      -- CP-element group 235: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Sample/$exit
      -- CP-element group 235: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Sample/ra
      -- 
    ra_5407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2057_inst_ack_0, ack => convolve_CP_4675_elements(235)); -- 
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	522 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	29 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_update_completed_
      -- CP-element group 236: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Update/$exit
      -- CP-element group 236: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2057_Update/ca
      -- 
    ca_5412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2057_inst_ack_1, ack => convolve_CP_4675_elements(236)); -- 
    -- CP-element group 237:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	160 
    -- CP-element group 237: 	176 
    -- CP-element group 237: 	144 
    -- CP-element group 237: marked-predecessors 
    -- CP-element group 237: 	239 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_sample_start_
      -- CP-element group 237: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Sample/$entry
      -- CP-element group 237: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Sample/rr
      -- 
    rr_5420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(237), ack => slice_2061_inst_req_0); -- 
    convolve_cp_element_group_237: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_237"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(239);
      gj_convolve_cp_element_group_237 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(237), clk => clk, reset => reset); --
    end block;
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	26 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: 	524 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_update_start_
      -- CP-element group 238: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Update/$entry
      -- CP-element group 238: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Update/cr
      -- 
    cr_5425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(238), ack => slice_2061_inst_req_1); -- 
    convolve_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(240) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: successors 
    -- CP-element group 239: marked-successors 
    -- CP-element group 239: 	158 
    -- CP-element group 239: 	174 
    -- CP-element group 239: 	142 
    -- CP-element group 239: 	237 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_sample_completed_
      -- CP-element group 239: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Sample/$exit
      -- CP-element group 239: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Sample/ra
      -- 
    ra_5421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 239_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2061_inst_ack_0, ack => convolve_CP_4675_elements(239)); -- 
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	522 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: 	29 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_update_completed_
      -- CP-element group 240: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Update/$exit
      -- CP-element group 240: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2061_Update/ca
      -- 
    ca_5426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2061_inst_ack_1, ack => convolve_CP_4675_elements(240)); -- 
    -- CP-element group 241:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	160 
    -- CP-element group 241: 	176 
    -- CP-element group 241: 	144 
    -- CP-element group 241: marked-predecessors 
    -- CP-element group 241: 	243 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	243 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_sample_start_
      -- CP-element group 241: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Sample/$entry
      -- CP-element group 241: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Sample/rr
      -- 
    rr_5434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(241), ack => slice_2065_inst_req_0); -- 
    convolve_cp_element_group_241: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_241"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(243);
      gj_convolve_cp_element_group_241 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(241), clk => clk, reset => reset); --
    end block;
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	26 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	524 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_update_start_
      -- CP-element group 242: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Update/$entry
      -- CP-element group 242: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Update/cr
      -- 
    cr_5439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(242), ack => slice_2065_inst_req_1); -- 
    convolve_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(244);
      gj_convolve_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	241 
    -- CP-element group 243: successors 
    -- CP-element group 243: marked-successors 
    -- CP-element group 243: 	158 
    -- CP-element group 243: 	174 
    -- CP-element group 243: 	142 
    -- CP-element group 243: 	241 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_sample_completed_
      -- CP-element group 243: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Sample/$exit
      -- CP-element group 243: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Sample/ra
      -- 
    ra_5435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2065_inst_ack_0, ack => convolve_CP_4675_elements(243)); -- 
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	522 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	29 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_update_completed_
      -- CP-element group 244: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Update/$exit
      -- CP-element group 244: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2065_Update/ca
      -- 
    ca_5440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2065_inst_ack_1, ack => convolve_CP_4675_elements(244)); -- 
    -- CP-element group 245:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	160 
    -- CP-element group 245: 	176 
    -- CP-element group 245: 	144 
    -- CP-element group 245: marked-predecessors 
    -- CP-element group 245: 	247 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	247 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_sample_start_
      -- CP-element group 245: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Sample/$entry
      -- CP-element group 245: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Sample/rr
      -- 
    rr_5448_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5448_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(245), ack => slice_2069_inst_req_0); -- 
    convolve_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(160) & convolve_CP_4675_elements(176) & convolve_CP_4675_elements(144) & convolve_CP_4675_elements(247);
      gj_convolve_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	26 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: 	524 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_update_start_
      -- CP-element group 246: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Update/$entry
      -- CP-element group 246: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Update/cr
      -- 
    cr_5453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(246), ack => slice_2069_inst_req_1); -- 
    convolve_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(248) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	245 
    -- CP-element group 247: successors 
    -- CP-element group 247: marked-successors 
    -- CP-element group 247: 	158 
    -- CP-element group 247: 	174 
    -- CP-element group 247: 	142 
    -- CP-element group 247: 	245 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_sample_completed_
      -- CP-element group 247: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Sample/$exit
      -- CP-element group 247: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Sample/ra
      -- 
    ra_5449_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2069_inst_ack_0, ack => convolve_CP_4675_elements(247)); -- 
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	522 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: 	29 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_update_completed_
      -- CP-element group 248: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Update/$exit
      -- CP-element group 248: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2069_Update/ca
      -- 
    ca_5454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2069_inst_ack_1, ack => convolve_CP_4675_elements(248)); -- 
    -- CP-element group 249:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	164 
    -- CP-element group 249: 	180 
    -- CP-element group 249: 	148 
    -- CP-element group 249: marked-predecessors 
    -- CP-element group 249: 	251 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	251 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Sample/rr
      -- 
    rr_5462_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5462_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(249), ack => slice_2073_inst_req_0); -- 
    convolve_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(251);
      gj_convolve_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	26 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: 	524 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_update_start_
      -- CP-element group 250: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Update/$entry
      -- CP-element group 250: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Update/cr
      -- 
    cr_5467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(250), ack => slice_2073_inst_req_1); -- 
    convolve_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(252) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	249 
    -- CP-element group 251: successors 
    -- CP-element group 251: marked-successors 
    -- CP-element group 251: 	162 
    -- CP-element group 251: 	249 
    -- CP-element group 251: 	146 
    -- CP-element group 251: 	178 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_sample_completed_
      -- CP-element group 251: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Sample/$exit
      -- CP-element group 251: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Sample/ra
      -- 
    ra_5463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2073_inst_ack_0, ack => convolve_CP_4675_elements(251)); -- 
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	522 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	48 
    -- CP-element group 252: 	29 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_update_completed_
      -- CP-element group 252: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Update/$exit
      -- CP-element group 252: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2073_Update/ca
      -- 
    ca_5468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2073_inst_ack_1, ack => convolve_CP_4675_elements(252)); -- 
    -- CP-element group 253:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	164 
    -- CP-element group 253: 	180 
    -- CP-element group 253: 	148 
    -- CP-element group 253: marked-predecessors 
    -- CP-element group 253: 	255 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	255 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_sample_start_
      -- CP-element group 253: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Sample/rr
      -- 
    rr_5476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(253), ack => slice_2077_inst_req_0); -- 
    convolve_cp_element_group_253: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_253"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(255);
      gj_convolve_cp_element_group_253 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(253), clk => clk, reset => reset); --
    end block;
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	26 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: 	524 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_update_start_
      -- CP-element group 254: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Update/$entry
      -- CP-element group 254: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Update/cr
      -- 
    cr_5481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(254), ack => slice_2077_inst_req_1); -- 
    convolve_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(256) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	253 
    -- CP-element group 255: successors 
    -- CP-element group 255: marked-successors 
    -- CP-element group 255: 	162 
    -- CP-element group 255: 	253 
    -- CP-element group 255: 	146 
    -- CP-element group 255: 	178 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_sample_completed_
      -- CP-element group 255: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Sample/$exit
      -- CP-element group 255: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Sample/ra
      -- 
    ra_5477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2077_inst_ack_0, ack => convolve_CP_4675_elements(255)); -- 
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	522 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	48 
    -- CP-element group 256: 	29 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_update_completed_
      -- CP-element group 256: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Update/$exit
      -- CP-element group 256: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2077_Update/ca
      -- 
    ca_5482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2077_inst_ack_1, ack => convolve_CP_4675_elements(256)); -- 
    -- CP-element group 257:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	164 
    -- CP-element group 257: 	180 
    -- CP-element group 257: 	148 
    -- CP-element group 257: marked-predecessors 
    -- CP-element group 257: 	259 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_sample_start_
      -- CP-element group 257: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Sample/$entry
      -- CP-element group 257: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Sample/rr
      -- 
    rr_5490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(257), ack => slice_2081_inst_req_0); -- 
    convolve_cp_element_group_257: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_257"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(259);
      gj_convolve_cp_element_group_257 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(257), clk => clk, reset => reset); --
    end block;
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	26 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: 	524 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_update_start_
      -- CP-element group 258: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Update/$entry
      -- CP-element group 258: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Update/cr
      -- 
    cr_5495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(258), ack => slice_2081_inst_req_1); -- 
    convolve_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(260) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: successors 
    -- CP-element group 259: marked-successors 
    -- CP-element group 259: 	162 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	146 
    -- CP-element group 259: 	178 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_sample_completed_
      -- CP-element group 259: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Sample/$exit
      -- CP-element group 259: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Sample/ra
      -- 
    ra_5491_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 259_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2081_inst_ack_0, ack => convolve_CP_4675_elements(259)); -- 
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	522 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	48 
    -- CP-element group 260: 	29 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_update_completed_
      -- CP-element group 260: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Update/$exit
      -- CP-element group 260: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2081_Update/ca
      -- 
    ca_5496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2081_inst_ack_1, ack => convolve_CP_4675_elements(260)); -- 
    -- CP-element group 261:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	164 
    -- CP-element group 261: 	180 
    -- CP-element group 261: 	148 
    -- CP-element group 261: marked-predecessors 
    -- CP-element group 261: 	263 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	263 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Sample/rr
      -- 
    rr_5504_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5504_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(261), ack => slice_2085_inst_req_0); -- 
    convolve_cp_element_group_261: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_261"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(263);
      gj_convolve_cp_element_group_261 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(261), clk => clk, reset => reset); --
    end block;
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	26 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	524 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_update_start_
      -- CP-element group 262: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Update/$entry
      -- CP-element group 262: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Update/cr
      -- 
    cr_5509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(262), ack => slice_2085_inst_req_1); -- 
    convolve_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(264);
      gj_convolve_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	261 
    -- CP-element group 263: successors 
    -- CP-element group 263: marked-successors 
    -- CP-element group 263: 	162 
    -- CP-element group 263: 	146 
    -- CP-element group 263: 	261 
    -- CP-element group 263: 	178 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_sample_completed_
      -- CP-element group 263: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Sample/$exit
      -- CP-element group 263: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Sample/ra
      -- 
    ra_5505_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2085_inst_ack_0, ack => convolve_CP_4675_elements(263)); -- 
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	522 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	48 
    -- CP-element group 264: 	29 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_update_completed_
      -- CP-element group 264: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Update/$exit
      -- CP-element group 264: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2085_Update/ca
      -- 
    ca_5510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2085_inst_ack_1, ack => convolve_CP_4675_elements(264)); -- 
    -- CP-element group 265:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	164 
    -- CP-element group 265: 	180 
    -- CP-element group 265: 	148 
    -- CP-element group 265: marked-predecessors 
    -- CP-element group 265: 	267 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	267 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Sample/rr
      -- CP-element group 265: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Sample/$entry
      -- CP-element group 265: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_sample_start_
      -- 
    rr_5518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(265), ack => slice_2089_inst_req_0); -- 
    convolve_cp_element_group_265: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_265"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(267);
      gj_convolve_cp_element_group_265 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(265), clk => clk, reset => reset); --
    end block;
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	26 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: 	524 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Update/$entry
      -- CP-element group 266: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Update/cr
      -- CP-element group 266: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_update_start_
      -- 
    cr_5523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(266), ack => slice_2089_inst_req_1); -- 
    convolve_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(268) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	265 
    -- CP-element group 267: successors 
    -- CP-element group 267: marked-successors 
    -- CP-element group 267: 	162 
    -- CP-element group 267: 	146 
    -- CP-element group 267: 	265 
    -- CP-element group 267: 	178 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Sample/ra
      -- CP-element group 267: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Sample/$exit
      -- CP-element group 267: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_sample_completed_
      -- 
    ra_5519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2089_inst_ack_0, ack => convolve_CP_4675_elements(267)); -- 
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	522 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	48 
    -- CP-element group 268: 	29 
    -- CP-element group 268: 	266 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Update/$exit
      -- CP-element group 268: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_Update/ca
      -- CP-element group 268: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2089_update_completed_
      -- 
    ca_5524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2089_inst_ack_1, ack => convolve_CP_4675_elements(268)); -- 
    -- CP-element group 269:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	164 
    -- CP-element group 269: 	180 
    -- CP-element group 269: 	148 
    -- CP-element group 269: marked-predecessors 
    -- CP-element group 269: 	271 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	271 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Sample/rr
      -- CP-element group 269: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_sample_start_
      -- CP-element group 269: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Sample/$entry
      -- 
    rr_5532_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5532_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(269), ack => slice_2093_inst_req_0); -- 
    convolve_cp_element_group_269: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_269"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(271);
      gj_convolve_cp_element_group_269 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(269), clk => clk, reset => reset); --
    end block;
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	26 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: 	524 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Update/$entry
      -- CP-element group 270: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Update/cr
      -- CP-element group 270: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_update_start_
      -- 
    cr_5537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(270), ack => slice_2093_inst_req_1); -- 
    convolve_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(272) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	269 
    -- CP-element group 271: successors 
    -- CP-element group 271: marked-successors 
    -- CP-element group 271: 	162 
    -- CP-element group 271: 	269 
    -- CP-element group 271: 	146 
    -- CP-element group 271: 	178 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Sample/ra
      -- CP-element group 271: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_sample_completed_
      -- CP-element group 271: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Sample/$exit
      -- 
    ra_5533_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2093_inst_ack_0, ack => convolve_CP_4675_elements(271)); -- 
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	522 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	48 
    -- CP-element group 272: 	29 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Update/$exit
      -- CP-element group 272: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_Update/ca
      -- CP-element group 272: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2093_update_completed_
      -- 
    ca_5538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2093_inst_ack_1, ack => convolve_CP_4675_elements(272)); -- 
    -- CP-element group 273:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	164 
    -- CP-element group 273: 	180 
    -- CP-element group 273: 	148 
    -- CP-element group 273: marked-predecessors 
    -- CP-element group 273: 	275 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	275 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Sample/$entry
      -- CP-element group 273: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Sample/rr
      -- CP-element group 273: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_sample_start_
      -- 
    rr_5546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(273), ack => slice_2097_inst_req_0); -- 
    convolve_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(275);
      gj_convolve_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	26 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: 	524 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Update/$entry
      -- CP-element group 274: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Update/cr
      -- CP-element group 274: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_update_start_
      -- 
    cr_5551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(274), ack => slice_2097_inst_req_1); -- 
    convolve_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(276) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	273 
    -- CP-element group 275: successors 
    -- CP-element group 275: marked-successors 
    -- CP-element group 275: 	162 
    -- CP-element group 275: 	273 
    -- CP-element group 275: 	146 
    -- CP-element group 275: 	178 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Sample/$exit
      -- CP-element group 275: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Sample/ra
      -- CP-element group 275: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_sample_completed_
      -- 
    ra_5547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2097_inst_ack_0, ack => convolve_CP_4675_elements(275)); -- 
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	522 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	48 
    -- CP-element group 276: 	29 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Update/$exit
      -- CP-element group 276: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_Update/ca
      -- CP-element group 276: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2097_update_completed_
      -- 
    ca_5552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2097_inst_ack_1, ack => convolve_CP_4675_elements(276)); -- 
    -- CP-element group 277:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	164 
    -- CP-element group 277: 	180 
    -- CP-element group 277: 	148 
    -- CP-element group 277: marked-predecessors 
    -- CP-element group 277: 	279 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_sample_start_
      -- CP-element group 277: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Sample/rr
      -- CP-element group 277: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Sample/$entry
      -- 
    rr_5560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(277), ack => slice_2101_inst_req_0); -- 
    convolve_cp_element_group_277: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_277"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(164) & convolve_CP_4675_elements(180) & convolve_CP_4675_elements(148) & convolve_CP_4675_elements(279);
      gj_convolve_cp_element_group_277 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(277), clk => clk, reset => reset); --
    end block;
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	26 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: 	524 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_update_start_
      -- CP-element group 278: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Update/$entry
      -- CP-element group 278: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Update/cr
      -- 
    cr_5565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(278), ack => slice_2101_inst_req_1); -- 
    convolve_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(280) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: successors 
    -- CP-element group 279: marked-successors 
    -- CP-element group 279: 	162 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	146 
    -- CP-element group 279: 	178 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Sample/$exit
      -- CP-element group 279: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Sample/ra
      -- CP-element group 279: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_sample_completed_
      -- 
    ra_5561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 279_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2101_inst_ack_0, ack => convolve_CP_4675_elements(279)); -- 
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	522 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: 	48 
    -- CP-element group 280: 	29 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_update_completed_
      -- CP-element group 280: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Update/$exit
      -- CP-element group 280: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2101_Update/ca
      -- 
    ca_5566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2101_inst_ack_1, ack => convolve_CP_4675_elements(280)); -- 
    -- CP-element group 281:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	184 
    -- CP-element group 281: 	168 
    -- CP-element group 281: 	152 
    -- CP-element group 281: marked-predecessors 
    -- CP-element group 281: 	283 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Sample/rr
      -- CP-element group 281: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Sample/$entry
      -- CP-element group 281: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_sample_start_
      -- 
    rr_5574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(281), ack => slice_2105_inst_req_0); -- 
    convolve_cp_element_group_281: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_281"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(283);
      gj_convolve_cp_element_group_281 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(281), clk => clk, reset => reset); --
    end block;
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	26 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: 	524 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_update_start_
      -- CP-element group 282: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Update/cr
      -- CP-element group 282: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Update/$entry
      -- 
    cr_5579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(282), ack => slice_2105_inst_req_1); -- 
    convolve_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(284) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: marked-successors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: 	182 
    -- CP-element group 283: 	166 
    -- CP-element group 283: 	150 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Sample/$exit
      -- CP-element group 283: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Sample/ra
      -- CP-element group 283: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_sample_completed_
      -- 
    ra_5575_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2105_inst_ack_0, ack => convolve_CP_4675_elements(283)); -- 
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	522 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	48 
    -- CP-element group 284: 	29 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_update_completed_
      -- CP-element group 284: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Update/ca
      -- CP-element group 284: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2105_Update/$exit
      -- 
    ca_5580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2105_inst_ack_1, ack => convolve_CP_4675_elements(284)); -- 
    -- CP-element group 285:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	184 
    -- CP-element group 285: 	168 
    -- CP-element group 285: 	152 
    -- CP-element group 285: marked-predecessors 
    -- CP-element group 285: 	287 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_sample_start_
      -- CP-element group 285: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Sample/$entry
      -- CP-element group 285: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Sample/rr
      -- 
    rr_5588_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5588_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(285), ack => slice_2109_inst_req_0); -- 
    convolve_cp_element_group_285: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_285"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(287);
      gj_convolve_cp_element_group_285 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(285), clk => clk, reset => reset); --
    end block;
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	26 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: 	524 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_update_start_
      -- CP-element group 286: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Update/$entry
      -- CP-element group 286: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Update/cr
      -- 
    cr_5593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(286), ack => slice_2109_inst_req_1); -- 
    convolve_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(288) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: successors 
    -- CP-element group 287: marked-successors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	182 
    -- CP-element group 287: 	166 
    -- CP-element group 287: 	150 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_sample_completed_
      -- CP-element group 287: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Sample/$exit
      -- CP-element group 287: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Sample/ra
      -- 
    ra_5589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 287_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2109_inst_ack_0, ack => convolve_CP_4675_elements(287)); -- 
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	522 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: 	48 
    -- CP-element group 288: 	29 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_update_completed_
      -- CP-element group 288: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Update/ca
      -- CP-element group 288: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2109_Update/$exit
      -- 
    ca_5594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2109_inst_ack_1, ack => convolve_CP_4675_elements(288)); -- 
    -- CP-element group 289:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	184 
    -- CP-element group 289: 	168 
    -- CP-element group 289: 	152 
    -- CP-element group 289: marked-predecessors 
    -- CP-element group 289: 	291 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	291 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Sample/$entry
      -- CP-element group 289: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Sample/rr
      -- CP-element group 289: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_sample_start_
      -- 
    rr_5602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(289), ack => slice_2113_inst_req_0); -- 
    convolve_cp_element_group_289: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_289"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(291);
      gj_convolve_cp_element_group_289 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(289), clk => clk, reset => reset); --
    end block;
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	26 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: 	524 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_update_start_
      -- CP-element group 290: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Update/$entry
      -- CP-element group 290: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Update/cr
      -- 
    cr_5607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(290), ack => slice_2113_inst_req_1); -- 
    convolve_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(292) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: successors 
    -- CP-element group 291: marked-successors 
    -- CP-element group 291: 	289 
    -- CP-element group 291: 	182 
    -- CP-element group 291: 	166 
    -- CP-element group 291: 	150 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Sample/ra
      -- CP-element group 291: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_sample_completed_
      -- 
    ra_5603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2113_inst_ack_0, ack => convolve_CP_4675_elements(291)); -- 
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	522 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: 	48 
    -- CP-element group 292: 	29 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_update_completed_
      -- CP-element group 292: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2113_Update/ca
      -- 
    ca_5608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2113_inst_ack_1, ack => convolve_CP_4675_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	184 
    -- CP-element group 293: 	168 
    -- CP-element group 293: 	152 
    -- CP-element group 293: marked-predecessors 
    -- CP-element group 293: 	295 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	295 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_sample_start_
      -- CP-element group 293: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Sample/$entry
      -- CP-element group 293: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Sample/rr
      -- 
    rr_5616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(293), ack => slice_2117_inst_req_0); -- 
    convolve_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(295);
      gj_convolve_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	26 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: 	524 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Update/cr
      -- CP-element group 294: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_update_start_
      -- CP-element group 294: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Update/$entry
      -- 
    cr_5621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(294), ack => slice_2117_inst_req_1); -- 
    convolve_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(296) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: successors 
    -- CP-element group 295: marked-successors 
    -- CP-element group 295: 	293 
    -- CP-element group 295: 	182 
    -- CP-element group 295: 	166 
    -- CP-element group 295: 	150 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_sample_completed_
      -- CP-element group 295: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Sample/$exit
      -- CP-element group 295: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Sample/ra
      -- 
    ra_5617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2117_inst_ack_0, ack => convolve_CP_4675_elements(295)); -- 
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	522 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: 	48 
    -- CP-element group 296: 	29 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Update/$exit
      -- CP-element group 296: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_update_completed_
      -- CP-element group 296: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2117_Update/ca
      -- 
    ca_5622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2117_inst_ack_1, ack => convolve_CP_4675_elements(296)); -- 
    -- CP-element group 297:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	184 
    -- CP-element group 297: 	168 
    -- CP-element group 297: 	152 
    -- CP-element group 297: marked-predecessors 
    -- CP-element group 297: 	299 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Sample/$entry
      -- CP-element group 297: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_sample_start_
      -- CP-element group 297: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Sample/rr
      -- 
    rr_5630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(297), ack => slice_2121_inst_req_0); -- 
    convolve_cp_element_group_297: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_297"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(299);
      gj_convolve_cp_element_group_297 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(297), clk => clk, reset => reset); --
    end block;
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	26 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: 	524 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_update_start_
      -- CP-element group 298: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Update/$entry
      -- CP-element group 298: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Update/cr
      -- 
    cr_5635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(298), ack => slice_2121_inst_req_1); -- 
    convolve_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(300) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: successors 
    -- CP-element group 299: marked-successors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: 	182 
    -- CP-element group 299: 	166 
    -- CP-element group 299: 	150 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_sample_completed_
      -- CP-element group 299: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Sample/$exit
      -- CP-element group 299: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Sample/ra
      -- 
    ra_5631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 299_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2121_inst_ack_0, ack => convolve_CP_4675_elements(299)); -- 
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	522 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	48 
    -- CP-element group 300: 	29 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_update_completed_
      -- CP-element group 300: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Update/$exit
      -- CP-element group 300: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2121_Update/ca
      -- 
    ca_5636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2121_inst_ack_1, ack => convolve_CP_4675_elements(300)); -- 
    -- CP-element group 301:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	184 
    -- CP-element group 301: 	168 
    -- CP-element group 301: 	152 
    -- CP-element group 301: marked-predecessors 
    -- CP-element group 301: 	303 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	303 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_sample_start_
      -- 
    rr_5644_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5644_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(301), ack => slice_2125_inst_req_0); -- 
    convolve_cp_element_group_301: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_301"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(303);
      gj_convolve_cp_element_group_301 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(301), clk => clk, reset => reset); --
    end block;
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	26 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: 	524 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_update_start_
      -- CP-element group 302: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Update/cr
      -- CP-element group 302: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Update/$entry
      -- 
    cr_5649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(302), ack => slice_2125_inst_req_1); -- 
    convolve_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(304) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: successors 
    -- CP-element group 303: marked-successors 
    -- CP-element group 303: 	301 
    -- CP-element group 303: 	182 
    -- CP-element group 303: 	166 
    -- CP-element group 303: 	150 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_sample_completed_
      -- CP-element group 303: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Sample/$exit
      -- CP-element group 303: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Sample/ra
      -- 
    ra_5645_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 303_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2125_inst_ack_0, ack => convolve_CP_4675_elements(303)); -- 
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	522 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	48 
    -- CP-element group 304: 	302 
    -- CP-element group 304: 	29 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Update/$exit
      -- CP-element group 304: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_Update/ca
      -- CP-element group 304: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2125_update_completed_
      -- 
    ca_5650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2125_inst_ack_1, ack => convolve_CP_4675_elements(304)); -- 
    -- CP-element group 305:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	184 
    -- CP-element group 305: 	168 
    -- CP-element group 305: 	152 
    -- CP-element group 305: marked-predecessors 
    -- CP-element group 305: 	307 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Sample/$entry
      -- CP-element group 305: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_sample_start_
      -- CP-element group 305: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Sample/rr
      -- 
    rr_5658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(305), ack => slice_2129_inst_req_0); -- 
    convolve_cp_element_group_305: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_305"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(307);
      gj_convolve_cp_element_group_305 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(305), clk => clk, reset => reset); --
    end block;
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	26 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: 	524 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Update/$entry
      -- CP-element group 306: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Update/cr
      -- CP-element group 306: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_update_start_
      -- 
    cr_5663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(306), ack => slice_2129_inst_req_1); -- 
    convolve_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(308) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: successors 
    -- CP-element group 307: marked-successors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	182 
    -- CP-element group 307: 	166 
    -- CP-element group 307: 	150 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Sample/ra
      -- CP-element group 307: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Sample/$exit
      -- CP-element group 307: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_sample_completed_
      -- 
    ra_5659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 307_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2129_inst_ack_0, ack => convolve_CP_4675_elements(307)); -- 
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	522 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: 	48 
    -- CP-element group 308: 	29 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Update/$exit
      -- CP-element group 308: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_Update/ca
      -- CP-element group 308: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2129_update_completed_
      -- 
    ca_5664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2129_inst_ack_1, ack => convolve_CP_4675_elements(308)); -- 
    -- CP-element group 309:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	184 
    -- CP-element group 309: 	168 
    -- CP-element group 309: 	152 
    -- CP-element group 309: marked-predecessors 
    -- CP-element group 309: 	311 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	311 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_sample_start_
      -- CP-element group 309: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Sample/rr
      -- 
    rr_5672_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5672_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(309), ack => slice_2133_inst_req_0); -- 
    convolve_cp_element_group_309: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_309"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(184) & convolve_CP_4675_elements(168) & convolve_CP_4675_elements(152) & convolve_CP_4675_elements(311);
      gj_convolve_cp_element_group_309 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(309), clk => clk, reset => reset); --
    end block;
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	26 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: 	524 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_update_start_
      -- CP-element group 310: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Update/cr
      -- 
    cr_5677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(310), ack => slice_2133_inst_req_1); -- 
    convolve_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(312) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: successors 
    -- CP-element group 311: marked-successors 
    -- CP-element group 311: 	309 
    -- CP-element group 311: 	182 
    -- CP-element group 311: 	166 
    -- CP-element group 311: 	150 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_sample_completed_
      -- CP-element group 311: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Sample/$exit
      -- CP-element group 311: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Sample/ra
      -- 
    ra_5673_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 311_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2133_inst_ack_0, ack => convolve_CP_4675_elements(311)); -- 
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: 	522 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: 	48 
    -- CP-element group 312: 	29 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_update_completed_
      -- CP-element group 312: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Update/$exit
      -- CP-element group 312: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2133_Update/ca
      -- 
    ca_5678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2133_inst_ack_1, ack => convolve_CP_4675_elements(312)); -- 
    -- CP-element group 313:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	156 
    -- CP-element group 313: 	172 
    -- CP-element group 313: 	188 
    -- CP-element group 313: marked-predecessors 
    -- CP-element group 313: 	315 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	315 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_sample_start_
      -- CP-element group 313: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Sample/$entry
      -- CP-element group 313: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Sample/rr
      -- 
    rr_5686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(313), ack => slice_2137_inst_req_0); -- 
    convolve_cp_element_group_313: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_313"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(315);
      gj_convolve_cp_element_group_313 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(313), clk => clk, reset => reset); --
    end block;
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	26 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: 	524 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_update_start_
      -- CP-element group 314: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Update/$entry
      -- CP-element group 314: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Update/cr
      -- 
    cr_5691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(314), ack => slice_2137_inst_req_1); -- 
    convolve_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(316) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: 	313 
    -- CP-element group 315: successors 
    -- CP-element group 315: marked-successors 
    -- CP-element group 315: 	154 
    -- CP-element group 315: 	313 
    -- CP-element group 315: 	186 
    -- CP-element group 315: 	170 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_sample_completed_
      -- CP-element group 315: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Sample/$exit
      -- CP-element group 315: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Sample/ra
      -- 
    ra_5687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 315_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2137_inst_ack_0, ack => convolve_CP_4675_elements(315)); -- 
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: 	522 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: 	48 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_update_completed_
      -- CP-element group 316: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Update/$exit
      -- CP-element group 316: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2137_Update/ca
      -- 
    ca_5692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2137_inst_ack_1, ack => convolve_CP_4675_elements(316)); -- 
    -- CP-element group 317:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	156 
    -- CP-element group 317: 	172 
    -- CP-element group 317: 	188 
    -- CP-element group 317: marked-predecessors 
    -- CP-element group 317: 	319 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	319 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_sample_start_
      -- CP-element group 317: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Sample/$entry
      -- CP-element group 317: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Sample/rr
      -- 
    rr_5700_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5700_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(317), ack => slice_2141_inst_req_0); -- 
    convolve_cp_element_group_317: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_317"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(319);
      gj_convolve_cp_element_group_317 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(317), clk => clk, reset => reset); --
    end block;
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	26 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: 	524 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_update_start_
      -- CP-element group 318: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Update/$entry
      -- CP-element group 318: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Update/cr
      -- 
    cr_5705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(318), ack => slice_2141_inst_req_1); -- 
    convolve_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(320) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: 	317 
    -- CP-element group 319: successors 
    -- CP-element group 319: marked-successors 
    -- CP-element group 319: 	154 
    -- CP-element group 319: 	317 
    -- CP-element group 319: 	186 
    -- CP-element group 319: 	170 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_sample_completed_
      -- CP-element group 319: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Sample/$exit
      -- CP-element group 319: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Sample/ra
      -- 
    ra_5701_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 319_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2141_inst_ack_0, ack => convolve_CP_4675_elements(319)); -- 
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: 	522 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: 	48 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_update_completed_
      -- CP-element group 320: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Update/$exit
      -- CP-element group 320: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2141_Update/ca
      -- 
    ca_5706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2141_inst_ack_1, ack => convolve_CP_4675_elements(320)); -- 
    -- CP-element group 321:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	156 
    -- CP-element group 321: 	172 
    -- CP-element group 321: 	188 
    -- CP-element group 321: marked-predecessors 
    -- CP-element group 321: 	323 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	323 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_sample_start_
      -- CP-element group 321: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Sample/$entry
      -- CP-element group 321: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Sample/rr
      -- 
    rr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5714_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(321), ack => slice_2145_inst_req_0); -- 
    convolve_cp_element_group_321: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_321"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(323);
      gj_convolve_cp_element_group_321 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(321), clk => clk, reset => reset); --
    end block;
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	26 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: 	524 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_update_start_
      -- CP-element group 322: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Update/$entry
      -- CP-element group 322: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Update/cr
      -- 
    cr_5719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(322), ack => slice_2145_inst_req_1); -- 
    convolve_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(324) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: 	321 
    -- CP-element group 323: successors 
    -- CP-element group 323: marked-successors 
    -- CP-element group 323: 	154 
    -- CP-element group 323: 	321 
    -- CP-element group 323: 	186 
    -- CP-element group 323: 	170 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_sample_completed_
      -- CP-element group 323: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Sample/$exit
      -- CP-element group 323: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Sample/ra
      -- 
    ra_5715_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 323_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2145_inst_ack_0, ack => convolve_CP_4675_elements(323)); -- 
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: 	522 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	48 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_update_completed_
      -- CP-element group 324: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Update/$exit
      -- CP-element group 324: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2145_Update/ca
      -- 
    ca_5720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2145_inst_ack_1, ack => convolve_CP_4675_elements(324)); -- 
    -- CP-element group 325:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	156 
    -- CP-element group 325: 	172 
    -- CP-element group 325: 	188 
    -- CP-element group 325: marked-predecessors 
    -- CP-element group 325: 	327 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	327 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_sample_start_
      -- CP-element group 325: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Sample/$entry
      -- CP-element group 325: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Sample/rr
      -- 
    rr_5728_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5728_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(325), ack => slice_2149_inst_req_0); -- 
    convolve_cp_element_group_325: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_325"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(327);
      gj_convolve_cp_element_group_325 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(325), clk => clk, reset => reset); --
    end block;
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	26 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: 	524 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_update_start_
      -- CP-element group 326: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Update/$entry
      -- CP-element group 326: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Update/cr
      -- 
    cr_5733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(326), ack => slice_2149_inst_req_1); -- 
    convolve_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(328) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: 	325 
    -- CP-element group 327: successors 
    -- CP-element group 327: marked-successors 
    -- CP-element group 327: 	154 
    -- CP-element group 327: 	325 
    -- CP-element group 327: 	186 
    -- CP-element group 327: 	170 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_sample_completed_
      -- CP-element group 327: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Sample/$exit
      -- CP-element group 327: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Sample/ra
      -- 
    ra_5729_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 327_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2149_inst_ack_0, ack => convolve_CP_4675_elements(327)); -- 
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: 	522 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: 	48 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_update_completed_
      -- CP-element group 328: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Update/$exit
      -- CP-element group 328: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2149_Update/ca
      -- 
    ca_5734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2149_inst_ack_1, ack => convolve_CP_4675_elements(328)); -- 
    -- CP-element group 329:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	156 
    -- CP-element group 329: 	172 
    -- CP-element group 329: 	188 
    -- CP-element group 329: marked-predecessors 
    -- CP-element group 329: 	331 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	331 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_sample_start_
      -- CP-element group 329: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Sample/$entry
      -- CP-element group 329: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Sample/rr
      -- 
    rr_5742_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5742_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(329), ack => slice_2153_inst_req_0); -- 
    convolve_cp_element_group_329: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_329"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(331);
      gj_convolve_cp_element_group_329 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(329), clk => clk, reset => reset); --
    end block;
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	26 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: 	524 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_update_start_
      -- CP-element group 330: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Update/$entry
      -- CP-element group 330: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Update/cr
      -- 
    cr_5747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(330), ack => slice_2153_inst_req_1); -- 
    convolve_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(332) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: 	329 
    -- CP-element group 331: successors 
    -- CP-element group 331: marked-successors 
    -- CP-element group 331: 	154 
    -- CP-element group 331: 	329 
    -- CP-element group 331: 	186 
    -- CP-element group 331: 	170 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_sample_completed_
      -- CP-element group 331: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Sample/$exit
      -- CP-element group 331: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Sample/ra
      -- 
    ra_5743_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 331_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2153_inst_ack_0, ack => convolve_CP_4675_elements(331)); -- 
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: 	522 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: 	48 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_update_completed_
      -- CP-element group 332: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Update/$exit
      -- CP-element group 332: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2153_Update/ca
      -- 
    ca_5748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2153_inst_ack_1, ack => convolve_CP_4675_elements(332)); -- 
    -- CP-element group 333:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	156 
    -- CP-element group 333: 	172 
    -- CP-element group 333: 	188 
    -- CP-element group 333: marked-predecessors 
    -- CP-element group 333: 	335 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	335 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_sample_start_
      -- CP-element group 333: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Sample/$entry
      -- CP-element group 333: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Sample/rr
      -- 
    rr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(333), ack => slice_2157_inst_req_0); -- 
    convolve_cp_element_group_333: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_333"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(335);
      gj_convolve_cp_element_group_333 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(333), clk => clk, reset => reset); --
    end block;
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	26 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: 	524 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_update_start_
      -- CP-element group 334: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Update/$entry
      -- CP-element group 334: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Update/cr
      -- 
    cr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(334), ack => slice_2157_inst_req_1); -- 
    convolve_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(336) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: 	333 
    -- CP-element group 335: successors 
    -- CP-element group 335: marked-successors 
    -- CP-element group 335: 	154 
    -- CP-element group 335: 	333 
    -- CP-element group 335: 	186 
    -- CP-element group 335: 	170 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_sample_completed_
      -- CP-element group 335: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Sample/$exit
      -- CP-element group 335: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Sample/ra
      -- 
    ra_5757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 335_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2157_inst_ack_0, ack => convolve_CP_4675_elements(335)); -- 
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: 	522 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: 	48 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_update_completed_
      -- CP-element group 336: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Update/$exit
      -- CP-element group 336: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2157_Update/ca
      -- 
    ca_5762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2157_inst_ack_1, ack => convolve_CP_4675_elements(336)); -- 
    -- CP-element group 337:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	156 
    -- CP-element group 337: 	172 
    -- CP-element group 337: 	188 
    -- CP-element group 337: marked-predecessors 
    -- CP-element group 337: 	339 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	339 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_sample_start_
      -- CP-element group 337: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Sample/$entry
      -- CP-element group 337: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Sample/rr
      -- 
    rr_5770_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5770_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(337), ack => slice_2161_inst_req_0); -- 
    convolve_cp_element_group_337: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_337"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(339);
      gj_convolve_cp_element_group_337 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(337), clk => clk, reset => reset); --
    end block;
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	26 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: 	524 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_update_start_
      -- CP-element group 338: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Update/$entry
      -- CP-element group 338: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Update/cr
      -- 
    cr_5775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(338), ack => slice_2161_inst_req_1); -- 
    convolve_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(340) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: 	337 
    -- CP-element group 339: successors 
    -- CP-element group 339: marked-successors 
    -- CP-element group 339: 	154 
    -- CP-element group 339: 	337 
    -- CP-element group 339: 	186 
    -- CP-element group 339: 	170 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_sample_completed_
      -- CP-element group 339: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Sample/$exit
      -- CP-element group 339: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Sample/ra
      -- 
    ra_5771_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 339_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2161_inst_ack_0, ack => convolve_CP_4675_elements(339)); -- 
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: 	522 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: 	48 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_update_completed_
      -- CP-element group 340: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Update/$exit
      -- CP-element group 340: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2161_Update/ca
      -- 
    ca_5776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2161_inst_ack_1, ack => convolve_CP_4675_elements(340)); -- 
    -- CP-element group 341:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	156 
    -- CP-element group 341: 	172 
    -- CP-element group 341: 	188 
    -- CP-element group 341: marked-predecessors 
    -- CP-element group 341: 	343 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	343 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_sample_start_
      -- CP-element group 341: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Sample/$entry
      -- CP-element group 341: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Sample/rr
      -- 
    rr_5784_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5784_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(341), ack => slice_2165_inst_req_0); -- 
    convolve_cp_element_group_341: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_341"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(156) & convolve_CP_4675_elements(172) & convolve_CP_4675_elements(188) & convolve_CP_4675_elements(343);
      gj_convolve_cp_element_group_341 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(341), clk => clk, reset => reset); --
    end block;
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	26 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: 	524 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_update_start_
      -- CP-element group 342: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Update/$entry
      -- CP-element group 342: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Update/cr
      -- 
    cr_5789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(342), ack => slice_2165_inst_req_1); -- 
    convolve_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(344) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: 	341 
    -- CP-element group 343: successors 
    -- CP-element group 343: marked-successors 
    -- CP-element group 343: 	154 
    -- CP-element group 343: 	341 
    -- CP-element group 343: 	186 
    -- CP-element group 343: 	170 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_sample_completed_
      -- CP-element group 343: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Sample/$exit
      -- CP-element group 343: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Sample/ra
      -- 
    ra_5785_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 343_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2165_inst_ack_0, ack => convolve_CP_4675_elements(343)); -- 
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: 	522 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: 	48 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_update_completed_
      -- CP-element group 344: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Update/$exit
      -- CP-element group 344: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2165_Update/ca
      -- 
    ca_5790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2165_inst_ack_1, ack => convolve_CP_4675_elements(344)); -- 
    -- CP-element group 345:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	23 
    -- CP-element group 345: marked-predecessors 
    -- CP-element group 345: 	348 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	347 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_sample_start_
      -- CP-element group 345: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Sample/$entry
      -- CP-element group 345: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Sample/rr
      -- 
    rr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5798_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(345), ack => RPIPE_kernel_pipe1_2306_inst_req_0); -- 
    convolve_cp_element_group_345: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_345"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(348);
      gj_convolve_cp_element_group_345 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(345), clk => clk, reset => reset); --
    end block;
    -- CP-element group 346:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	347 
    -- CP-element group 346: 	72 
    -- CP-element group 346: 	91 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	407 
    -- CP-element group 346: 	411 
    -- CP-element group 346: 	391 
    -- CP-element group 346: 	383 
    -- CP-element group 346: 	387 
    -- CP-element group 346: 	403 
    -- CP-element group 346: 	395 
    -- CP-element group 346: 	399 
    -- CP-element group 346: 	494 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: marked-successors 
    -- CP-element group 346: 	87 
    -- CP-element group 346: 	68 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_update_start_
      -- CP-element group 346: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Update/$entry
      -- CP-element group 346: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Update/cr
      -- 
    cr_5803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(346), ack => RPIPE_kernel_pipe1_2306_inst_req_1); -- 
    convolve_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 15,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(347) & convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(407) & convolve_CP_4675_elements(411) & convolve_CP_4675_elements(391) & convolve_CP_4675_elements(383) & convolve_CP_4675_elements(387) & convolve_CP_4675_elements(403) & convolve_CP_4675_elements(395) & convolve_CP_4675_elements(399) & convolve_CP_4675_elements(494);
      gj_convolve_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  transition  input  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: 	345 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	346 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_sample_completed_
      -- CP-element group 347: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Sample/$exit
      -- CP-element group 347: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Sample/ra
      -- 
    ra_5799_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 347_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2306_inst_ack_0, ack => convolve_CP_4675_elements(347)); -- 
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: 	409 
    -- CP-element group 348: 	389 
    -- CP-element group 348: 	393 
    -- CP-element group 348: 	381 
    -- CP-element group 348: 	385 
    -- CP-element group 348: 	401 
    -- CP-element group 348: 	405 
    -- CP-element group 348: 	397 
    -- CP-element group 348: 	493 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	345 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_update_completed_
      -- CP-element group 348: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Update/$exit
      -- CP-element group 348: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe1_2306_Update/ca
      -- 
    ca_5804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe1_2306_inst_ack_1, ack => convolve_CP_4675_elements(348)); -- 
    -- CP-element group 349:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	23 
    -- CP-element group 349: marked-predecessors 
    -- CP-element group 349: 	352 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	351 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_sample_start_
      -- CP-element group 349: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Sample/$entry
      -- CP-element group 349: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Sample/rr
      -- 
    rr_5812_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5812_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(349), ack => RPIPE_kernel_pipe2_2310_inst_req_0); -- 
    convolve_cp_element_group_349: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_349"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(352);
      gj_convolve_cp_element_group_349 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(349), clk => clk, reset => reset); --
    end block;
    -- CP-element group 350:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	72 
    -- CP-element group 350: 	351 
    -- CP-element group 350: 	91 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	419 
    -- CP-element group 350: 	423 
    -- CP-element group 350: 	439 
    -- CP-element group 350: 	443 
    -- CP-element group 350: 	427 
    -- CP-element group 350: 	501 
    -- CP-element group 350: 	415 
    -- CP-element group 350: 	431 
    -- CP-element group 350: 	435 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: marked-successors 
    -- CP-element group 350: 	87 
    -- CP-element group 350: 	68 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_update_start_
      -- CP-element group 350: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Update/$entry
      -- CP-element group 350: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Update/cr
      -- 
    cr_5817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(350), ack => RPIPE_kernel_pipe2_2310_inst_req_1); -- 
    convolve_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(351) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(419) & convolve_CP_4675_elements(423) & convolve_CP_4675_elements(439) & convolve_CP_4675_elements(443) & convolve_CP_4675_elements(427) & convolve_CP_4675_elements(501) & convolve_CP_4675_elements(415) & convolve_CP_4675_elements(431) & convolve_CP_4675_elements(435);
      gj_convolve_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  transition  input  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: 	349 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	350 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_sample_completed_
      -- CP-element group 351: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Sample/$exit
      -- CP-element group 351: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Sample/ra
      -- 
    ra_5813_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 351_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2310_inst_ack_0, ack => convolve_CP_4675_elements(351)); -- 
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: 	421 
    -- CP-element group 352: 	437 
    -- CP-element group 352: 	441 
    -- CP-element group 352: 	425 
    -- CP-element group 352: 	429 
    -- CP-element group 352: 	500 
    -- CP-element group 352: 	413 
    -- CP-element group 352: 	417 
    -- CP-element group 352: 	433 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	349 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_update_completed_
      -- CP-element group 352: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Update/$exit
      -- CP-element group 352: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe2_2310_Update/ca
      -- 
    ca_5818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe2_2310_inst_ack_1, ack => convolve_CP_4675_elements(352)); -- 
    -- CP-element group 353:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	23 
    -- CP-element group 353: marked-predecessors 
    -- CP-element group 353: 	356 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	355 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_sample_start_
      -- CP-element group 353: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Sample/$entry
      -- CP-element group 353: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Sample/rr
      -- 
    rr_5826_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5826_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(353), ack => RPIPE_kernel_pipe3_2314_inst_req_0); -- 
    convolve_cp_element_group_353: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_353"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(356);
      gj_convolve_cp_element_group_353 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(353), clk => clk, reset => reset); --
    end block;
    -- CP-element group 354:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	72 
    -- CP-element group 354: 	355 
    -- CP-element group 354: 	91 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	463 
    -- CP-element group 354: 	475 
    -- CP-element group 354: 	451 
    -- CP-element group 354: 	455 
    -- CP-element group 354: 	459 
    -- CP-element group 354: 	447 
    -- CP-element group 354: 	467 
    -- CP-element group 354: 	471 
    -- CP-element group 354: 	508 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: marked-successors 
    -- CP-element group 354: 	87 
    -- CP-element group 354: 	68 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_update_start_
      -- CP-element group 354: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Update/$entry
      -- CP-element group 354: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Update/cr
      -- 
    cr_5831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(354), ack => RPIPE_kernel_pipe3_2314_inst_req_1); -- 
    convolve_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(355) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(463) & convolve_CP_4675_elements(475) & convolve_CP_4675_elements(451) & convolve_CP_4675_elements(455) & convolve_CP_4675_elements(459) & convolve_CP_4675_elements(447) & convolve_CP_4675_elements(467) & convolve_CP_4675_elements(471) & convolve_CP_4675_elements(508);
      gj_convolve_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  transition  input  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: 	353 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	354 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_sample_completed_
      -- CP-element group 355: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Sample/$exit
      -- CP-element group 355: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Sample/ra
      -- 
    ra_5827_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 355_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2314_inst_ack_0, ack => convolve_CP_4675_elements(355)); -- 
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: 	461 
    -- CP-element group 356: 	465 
    -- CP-element group 356: 	473 
    -- CP-element group 356: 	449 
    -- CP-element group 356: 	453 
    -- CP-element group 356: 	457 
    -- CP-element group 356: 	445 
    -- CP-element group 356: 	469 
    -- CP-element group 356: 	507 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	353 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_update_completed_
      -- CP-element group 356: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Update/$exit
      -- CP-element group 356: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_kernel_pipe3_2314_Update/ca
      -- 
    ca_5832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_kernel_pipe3_2314_inst_ack_1, ack => convolve_CP_4675_elements(356)); -- 
    -- CP-element group 357:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	23 
    -- CP-element group 357: marked-predecessors 
    -- CP-element group 357: 	360 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	359 
    -- CP-element group 357:  members (3) 
      -- CP-element group 357: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_sample_start_
      -- CP-element group 357: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Sample/$entry
      -- CP-element group 357: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Sample/rr
      -- 
    rr_5840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(357), ack => RPIPE_xxconvolvexxconv_k1_2318_inst_req_0); -- 
    convolve_cp_element_group_357: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_357"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(360);
      gj_convolve_cp_element_group_357 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(357), clk => clk, reset => reset); --
    end block;
    -- CP-element group 358:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	72 
    -- CP-element group 358: 	359 
    -- CP-element group 358: 	91 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	407 
    -- CP-element group 358: 	411 
    -- CP-element group 358: 	391 
    -- CP-element group 358: 	383 
    -- CP-element group 358: 	387 
    -- CP-element group 358: 	403 
    -- CP-element group 358: 	395 
    -- CP-element group 358: 	399 
    -- CP-element group 358: 	494 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: marked-successors 
    -- CP-element group 358: 	87 
    -- CP-element group 358: 	68 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_update_start_
      -- CP-element group 358: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Update/$entry
      -- CP-element group 358: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Update/cr
      -- 
    cr_5845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(358), ack => RPIPE_xxconvolvexxconv_k1_2318_inst_req_1); -- 
    convolve_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 1,2 => 15,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(359) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(407) & convolve_CP_4675_elements(411) & convolve_CP_4675_elements(391) & convolve_CP_4675_elements(383) & convolve_CP_4675_elements(387) & convolve_CP_4675_elements(403) & convolve_CP_4675_elements(395) & convolve_CP_4675_elements(399) & convolve_CP_4675_elements(494);
      gj_convolve_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  transition  input  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: 	357 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	358 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_sample_completed_
      -- CP-element group 359: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Sample/$exit
      -- CP-element group 359: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Sample/ra
      -- 
    ra_5841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 359_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2318_inst_ack_0, ack => convolve_CP_4675_elements(359)); -- 
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: 	409 
    -- CP-element group 360: 	389 
    -- CP-element group 360: 	393 
    -- CP-element group 360: 	381 
    -- CP-element group 360: 	385 
    -- CP-element group 360: 	401 
    -- CP-element group 360: 	405 
    -- CP-element group 360: 	397 
    -- CP-element group 360: 	493 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	357 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_update_completed_
      -- CP-element group 360: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Update/$exit
      -- CP-element group 360: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k1_2318_Update/ca
      -- 
    ca_5846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k1_2318_inst_ack_1, ack => convolve_CP_4675_elements(360)); -- 
    -- CP-element group 361:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	23 
    -- CP-element group 361: marked-predecessors 
    -- CP-element group 361: 	364 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	363 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_sample_start_
      -- CP-element group 361: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Sample/$entry
      -- CP-element group 361: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Sample/rr
      -- 
    rr_5854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(361), ack => RPIPE_xxconvolvexxconv_k2_2322_inst_req_0); -- 
    convolve_cp_element_group_361: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_361"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(364);
      gj_convolve_cp_element_group_361 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(361), clk => clk, reset => reset); --
    end block;
    -- CP-element group 362:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	72 
    -- CP-element group 362: 	91 
    -- CP-element group 362: 	363 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	419 
    -- CP-element group 362: 	423 
    -- CP-element group 362: 	439 
    -- CP-element group 362: 	443 
    -- CP-element group 362: 	427 
    -- CP-element group 362: 	501 
    -- CP-element group 362: 	415 
    -- CP-element group 362: 	431 
    -- CP-element group 362: 	435 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: marked-successors 
    -- CP-element group 362: 	87 
    -- CP-element group 362: 	68 
    -- CP-element group 362:  members (3) 
      -- CP-element group 362: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_update_start_
      -- CP-element group 362: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Update/$entry
      -- CP-element group 362: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Update/cr
      -- 
    cr_5859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(362), ack => RPIPE_xxconvolvexxconv_k2_2322_inst_req_1); -- 
    convolve_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(363) & convolve_CP_4675_elements(419) & convolve_CP_4675_elements(423) & convolve_CP_4675_elements(439) & convolve_CP_4675_elements(443) & convolve_CP_4675_elements(427) & convolve_CP_4675_elements(501) & convolve_CP_4675_elements(415) & convolve_CP_4675_elements(431) & convolve_CP_4675_elements(435);
      gj_convolve_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  transition  input  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: 	361 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	362 
    -- CP-element group 363:  members (3) 
      -- CP-element group 363: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_sample_completed_
      -- CP-element group 363: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Sample/$exit
      -- CP-element group 363: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Sample/ra
      -- 
    ra_5855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 363_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2322_inst_ack_0, ack => convolve_CP_4675_elements(363)); -- 
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	421 
    -- CP-element group 364: 	437 
    -- CP-element group 364: 	441 
    -- CP-element group 364: 	425 
    -- CP-element group 364: 	429 
    -- CP-element group 364: 	500 
    -- CP-element group 364: 	413 
    -- CP-element group 364: 	417 
    -- CP-element group 364: 	433 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	361 
    -- CP-element group 364:  members (3) 
      -- CP-element group 364: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_update_completed_
      -- CP-element group 364: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Update/$exit
      -- CP-element group 364: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k2_2322_Update/ca
      -- 
    ca_5860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k2_2322_inst_ack_1, ack => convolve_CP_4675_elements(364)); -- 
    -- CP-element group 365:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	23 
    -- CP-element group 365: marked-predecessors 
    -- CP-element group 365: 	368 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	367 
    -- CP-element group 365:  members (3) 
      -- CP-element group 365: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_sample_start_
      -- CP-element group 365: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Sample/$entry
      -- CP-element group 365: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Sample/rr
      -- 
    rr_5868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(365), ack => RPIPE_xxconvolvexxconv_k3_2326_inst_req_0); -- 
    convolve_cp_element_group_365: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_365"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(368);
      gj_convolve_cp_element_group_365 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(365), clk => clk, reset => reset); --
    end block;
    -- CP-element group 366:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	72 
    -- CP-element group 366: 	91 
    -- CP-element group 366: 	367 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	463 
    -- CP-element group 366: 	475 
    -- CP-element group 366: 	451 
    -- CP-element group 366: 	455 
    -- CP-element group 366: 	459 
    -- CP-element group 366: 	447 
    -- CP-element group 366: 	467 
    -- CP-element group 366: 	471 
    -- CP-element group 366: 	508 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366: marked-successors 
    -- CP-element group 366: 	87 
    -- CP-element group 366: 	68 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_update_start_
      -- CP-element group 366: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Update/$entry
      -- CP-element group 366: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Update/cr
      -- 
    cr_5873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(366), ack => RPIPE_xxconvolvexxconv_k3_2326_inst_req_1); -- 
    convolve_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 15,1 => 15,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(367) & convolve_CP_4675_elements(463) & convolve_CP_4675_elements(475) & convolve_CP_4675_elements(451) & convolve_CP_4675_elements(455) & convolve_CP_4675_elements(459) & convolve_CP_4675_elements(447) & convolve_CP_4675_elements(467) & convolve_CP_4675_elements(471) & convolve_CP_4675_elements(508);
      gj_convolve_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  transition  input  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: 	365 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	366 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_sample_completed_
      -- CP-element group 367: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Sample/$exit
      -- CP-element group 367: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Sample/ra
      -- 
    ra_5869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 367_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2326_inst_ack_0, ack => convolve_CP_4675_elements(367)); -- 
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: successors 
    -- CP-element group 368: 	461 
    -- CP-element group 368: 	465 
    -- CP-element group 368: 	473 
    -- CP-element group 368: 	449 
    -- CP-element group 368: 	453 
    -- CP-element group 368: 	457 
    -- CP-element group 368: 	445 
    -- CP-element group 368: 	469 
    -- CP-element group 368: 	507 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	365 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_update_completed_
      -- CP-element group 368: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Update/$exit
      -- CP-element group 368: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/RPIPE_xxconvolvexxconv_k3_2326_Update/ca
      -- 
    ca_5874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_xxconvolvexxconv_k3_2326_inst_ack_1, ack => convolve_CP_4675_elements(368)); -- 
    -- CP-element group 369:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	72 
    -- CP-element group 369: 	91 
    -- CP-element group 369: marked-predecessors 
    -- CP-element group 369: 	371 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	371 
    -- CP-element group 369:  members (3) 
      -- CP-element group 369: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_sample_start_
      -- CP-element group 369: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Sample/$entry
      -- CP-element group 369: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Sample/req
      -- 
    req_5882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(369), ack => W_read_k_2284_delayed_1_0_2328_inst_req_0); -- 
    convolve_cp_element_group_369: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_369"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(371);
      gj_convolve_cp_element_group_369 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(369), clk => clk, reset => reset); --
    end block;
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	407 
    -- CP-element group 370: 	411 
    -- CP-element group 370: 	391 
    -- CP-element group 370: 	383 
    -- CP-element group 370: 	387 
    -- CP-element group 370: 	372 
    -- CP-element group 370: 	403 
    -- CP-element group 370: 	395 
    -- CP-element group 370: 	399 
    -- CP-element group 370: 	494 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_update_start_
      -- CP-element group 370: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Update/$entry
      -- CP-element group 370: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Update/req
      -- 
    req_5887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(370), ack => W_read_k_2284_delayed_1_0_2328_inst_req_1); -- 
    convolve_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(407) & convolve_CP_4675_elements(411) & convolve_CP_4675_elements(391) & convolve_CP_4675_elements(383) & convolve_CP_4675_elements(387) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(403) & convolve_CP_4675_elements(395) & convolve_CP_4675_elements(399) & convolve_CP_4675_elements(494);
      gj_convolve_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: successors 
    -- CP-element group 371: marked-successors 
    -- CP-element group 371: 	369 
    -- CP-element group 371: 	87 
    -- CP-element group 371: 	68 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_sample_completed_
      -- CP-element group 371: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Sample/$exit
      -- CP-element group 371: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Sample/ack
      -- 
    ack_5883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 371_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2284_delayed_1_0_2328_inst_ack_0, ack => convolve_CP_4675_elements(371)); -- 
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: successors 
    -- CP-element group 372: 	409 
    -- CP-element group 372: 	389 
    -- CP-element group 372: 	393 
    -- CP-element group 372: 	381 
    -- CP-element group 372: 	385 
    -- CP-element group 372: 	401 
    -- CP-element group 372: 	405 
    -- CP-element group 372: 	397 
    -- CP-element group 372: 	493 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_update_completed_
      -- CP-element group 372: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Update/$exit
      -- CP-element group 372: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2330_Update/ack
      -- 
    ack_5888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2284_delayed_1_0_2328_inst_ack_1, ack => convolve_CP_4675_elements(372)); -- 
    -- CP-element group 373:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	72 
    -- CP-element group 373: 	91 
    -- CP-element group 373: marked-predecessors 
    -- CP-element group 373: 	375 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	375 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_sample_start_
      -- CP-element group 373: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Sample/$entry
      -- CP-element group 373: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Sample/req
      -- 
    req_5896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(373), ack => W_read_k_2290_delayed_1_0_2337_inst_req_0); -- 
    convolve_cp_element_group_373: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_373"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(375);
      gj_convolve_cp_element_group_373 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(373), clk => clk, reset => reset); --
    end block;
    -- CP-element group 374:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: marked-predecessors 
    -- CP-element group 374: 	419 
    -- CP-element group 374: 	423 
    -- CP-element group 374: 	439 
    -- CP-element group 374: 	443 
    -- CP-element group 374: 	427 
    -- CP-element group 374: 	501 
    -- CP-element group 374: 	415 
    -- CP-element group 374: 	376 
    -- CP-element group 374: 	431 
    -- CP-element group 374: 	435 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (3) 
      -- CP-element group 374: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_update_start_
      -- CP-element group 374: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Update/$entry
      -- CP-element group 374: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Update/req
      -- 
    req_5901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(374), ack => W_read_k_2290_delayed_1_0_2337_inst_req_1); -- 
    convolve_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(419) & convolve_CP_4675_elements(423) & convolve_CP_4675_elements(439) & convolve_CP_4675_elements(443) & convolve_CP_4675_elements(427) & convolve_CP_4675_elements(501) & convolve_CP_4675_elements(415) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(431) & convolve_CP_4675_elements(435);
      gj_convolve_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: successors 
    -- CP-element group 375: marked-successors 
    -- CP-element group 375: 	373 
    -- CP-element group 375: 	87 
    -- CP-element group 375: 	68 
    -- CP-element group 375:  members (3) 
      -- CP-element group 375: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_sample_completed_
      -- CP-element group 375: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Sample/$exit
      -- CP-element group 375: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Sample/ack
      -- 
    ack_5897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 375_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2290_delayed_1_0_2337_inst_ack_0, ack => convolve_CP_4675_elements(375)); -- 
    -- CP-element group 376:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	421 
    -- CP-element group 376: 	437 
    -- CP-element group 376: 	441 
    -- CP-element group 376: 	425 
    -- CP-element group 376: 	429 
    -- CP-element group 376: 	500 
    -- CP-element group 376: 	413 
    -- CP-element group 376: 	417 
    -- CP-element group 376: 	433 
    -- CP-element group 376: marked-successors 
    -- CP-element group 376: 	374 
    -- CP-element group 376:  members (3) 
      -- CP-element group 376: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_update_completed_
      -- CP-element group 376: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Update/$exit
      -- CP-element group 376: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2339_Update/ack
      -- 
    ack_5902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2290_delayed_1_0_2337_inst_ack_1, ack => convolve_CP_4675_elements(376)); -- 
    -- CP-element group 377:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	72 
    -- CP-element group 377: 	91 
    -- CP-element group 377: marked-predecessors 
    -- CP-element group 377: 	379 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	379 
    -- CP-element group 377:  members (3) 
      -- CP-element group 377: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_sample_start_
      -- CP-element group 377: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Sample/$entry
      -- CP-element group 377: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Sample/req
      -- 
    req_5910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(377), ack => W_read_k_2296_delayed_1_0_2346_inst_req_0); -- 
    convolve_cp_element_group_377: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_377"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(379);
      gj_convolve_cp_element_group_377 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(377), clk => clk, reset => reset); --
    end block;
    -- CP-element group 378:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: marked-predecessors 
    -- CP-element group 378: 	463 
    -- CP-element group 378: 	475 
    -- CP-element group 378: 	451 
    -- CP-element group 378: 	455 
    -- CP-element group 378: 	459 
    -- CP-element group 378: 	447 
    -- CP-element group 378: 	467 
    -- CP-element group 378: 	471 
    -- CP-element group 378: 	508 
    -- CP-element group 378: 	380 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_update_start_
      -- CP-element group 378: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Update/$entry
      -- CP-element group 378: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Update/req
      -- 
    req_5915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(378), ack => W_read_k_2296_delayed_1_0_2346_inst_req_1); -- 
    convolve_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(463) & convolve_CP_4675_elements(475) & convolve_CP_4675_elements(451) & convolve_CP_4675_elements(455) & convolve_CP_4675_elements(459) & convolve_CP_4675_elements(447) & convolve_CP_4675_elements(467) & convolve_CP_4675_elements(471) & convolve_CP_4675_elements(508) & convolve_CP_4675_elements(380);
      gj_convolve_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: 	377 
    -- CP-element group 379: successors 
    -- CP-element group 379: marked-successors 
    -- CP-element group 379: 	87 
    -- CP-element group 379: 	68 
    -- CP-element group 379: 	377 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_sample_completed_
      -- CP-element group 379: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Sample/$exit
      -- CP-element group 379: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Sample/ack
      -- 
    ack_5911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 379_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2296_delayed_1_0_2346_inst_ack_0, ack => convolve_CP_4675_elements(379)); -- 
    -- CP-element group 380:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: 	461 
    -- CP-element group 380: 	465 
    -- CP-element group 380: 	473 
    -- CP-element group 380: 	449 
    -- CP-element group 380: 	453 
    -- CP-element group 380: 	457 
    -- CP-element group 380: 	445 
    -- CP-element group 380: 	469 
    -- CP-element group 380: 	507 
    -- CP-element group 380: marked-successors 
    -- CP-element group 380: 	378 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_update_completed_
      -- CP-element group 380: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Update/$exit
      -- CP-element group 380: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2348_Update/ack
      -- 
    ack_5916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_k_2296_delayed_1_0_2346_inst_ack_1, ack => convolve_CP_4675_elements(380)); -- 
    -- CP-element group 381:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	348 
    -- CP-element group 381: 	360 
    -- CP-element group 381: 	372 
    -- CP-element group 381: marked-predecessors 
    -- CP-element group 381: 	383 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	383 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_sample_start_
      -- CP-element group 381: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Sample/$entry
      -- CP-element group 381: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Sample/rr
      -- 
    rr_5924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(381), ack => slice_2357_inst_req_0); -- 
    convolve_cp_element_group_381: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_381"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(383);
      gj_convolve_cp_element_group_381 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(381), clk => clk, reset => reset); --
    end block;
    -- CP-element group 382:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	26 
    -- CP-element group 382: marked-predecessors 
    -- CP-element group 382: 	384 
    -- CP-element group 382: 	524 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	384 
    -- CP-element group 382:  members (3) 
      -- CP-element group 382: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_update_start_
      -- CP-element group 382: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Update/$entry
      -- CP-element group 382: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Update/cr
      -- 
    cr_5929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(382), ack => slice_2357_inst_req_1); -- 
    convolve_cp_element_group_382: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_382"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(384) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_382 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(382), clk => clk, reset => reset); --
    end block;
    -- CP-element group 383:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	381 
    -- CP-element group 383: successors 
    -- CP-element group 383: marked-successors 
    -- CP-element group 383: 	346 
    -- CP-element group 383: 	358 
    -- CP-element group 383: 	381 
    -- CP-element group 383: 	370 
    -- CP-element group 383:  members (3) 
      -- CP-element group 383: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_sample_completed_
      -- CP-element group 383: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Sample/$exit
      -- CP-element group 383: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Sample/ra
      -- 
    ra_5925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 383_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2357_inst_ack_0, ack => convolve_CP_4675_elements(383)); -- 
    -- CP-element group 384:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	522 
    -- CP-element group 384: marked-successors 
    -- CP-element group 384: 	382 
    -- CP-element group 384: 	48 
    -- CP-element group 384: 	29 
    -- CP-element group 384:  members (3) 
      -- CP-element group 384: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_update_completed_
      -- CP-element group 384: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Update/$exit
      -- CP-element group 384: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2357_Update/ca
      -- 
    ca_5930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 384_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2357_inst_ack_1, ack => convolve_CP_4675_elements(384)); -- 
    -- CP-element group 385:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	348 
    -- CP-element group 385: 	360 
    -- CP-element group 385: 	372 
    -- CP-element group 385: marked-predecessors 
    -- CP-element group 385: 	387 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	387 
    -- CP-element group 385:  members (3) 
      -- CP-element group 385: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_sample_start_
      -- CP-element group 385: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Sample/$entry
      -- CP-element group 385: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Sample/rr
      -- 
    rr_5938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(385), ack => slice_2361_inst_req_0); -- 
    convolve_cp_element_group_385: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_385"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(387);
      gj_convolve_cp_element_group_385 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(385), clk => clk, reset => reset); --
    end block;
    -- CP-element group 386:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	26 
    -- CP-element group 386: marked-predecessors 
    -- CP-element group 386: 	388 
    -- CP-element group 386: 	524 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	388 
    -- CP-element group 386:  members (3) 
      -- CP-element group 386: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_update_start_
      -- CP-element group 386: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Update/$entry
      -- CP-element group 386: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Update/cr
      -- 
    cr_5943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(386), ack => slice_2361_inst_req_1); -- 
    convolve_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(388) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	385 
    -- CP-element group 387: successors 
    -- CP-element group 387: marked-successors 
    -- CP-element group 387: 	346 
    -- CP-element group 387: 	358 
    -- CP-element group 387: 	385 
    -- CP-element group 387: 	370 
    -- CP-element group 387:  members (3) 
      -- CP-element group 387: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_sample_completed_
      -- CP-element group 387: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Sample/$exit
      -- CP-element group 387: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Sample/ra
      -- 
    ra_5939_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2361_inst_ack_0, ack => convolve_CP_4675_elements(387)); -- 
    -- CP-element group 388:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: successors 
    -- CP-element group 388: 	522 
    -- CP-element group 388: marked-successors 
    -- CP-element group 388: 	386 
    -- CP-element group 388: 	48 
    -- CP-element group 388: 	29 
    -- CP-element group 388:  members (3) 
      -- CP-element group 388: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_update_completed_
      -- CP-element group 388: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Update/$exit
      -- CP-element group 388: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2361_Update/ca
      -- 
    ca_5944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2361_inst_ack_1, ack => convolve_CP_4675_elements(388)); -- 
    -- CP-element group 389:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	348 
    -- CP-element group 389: 	360 
    -- CP-element group 389: 	372 
    -- CP-element group 389: marked-predecessors 
    -- CP-element group 389: 	391 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	391 
    -- CP-element group 389:  members (3) 
      -- CP-element group 389: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_sample_start_
      -- CP-element group 389: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Sample/$entry
      -- CP-element group 389: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Sample/rr
      -- 
    rr_5952_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5952_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(389), ack => slice_2365_inst_req_0); -- 
    convolve_cp_element_group_389: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_389"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(391);
      gj_convolve_cp_element_group_389 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(389), clk => clk, reset => reset); --
    end block;
    -- CP-element group 390:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	26 
    -- CP-element group 390: marked-predecessors 
    -- CP-element group 390: 	392 
    -- CP-element group 390: 	524 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	392 
    -- CP-element group 390:  members (3) 
      -- CP-element group 390: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_update_start_
      -- CP-element group 390: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Update/cr
      -- 
    cr_5957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(390), ack => slice_2365_inst_req_1); -- 
    convolve_cp_element_group_390: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_390"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(392) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_390 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(390), clk => clk, reset => reset); --
    end block;
    -- CP-element group 391:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	389 
    -- CP-element group 391: successors 
    -- CP-element group 391: marked-successors 
    -- CP-element group 391: 	346 
    -- CP-element group 391: 	358 
    -- CP-element group 391: 	389 
    -- CP-element group 391: 	370 
    -- CP-element group 391:  members (3) 
      -- CP-element group 391: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_sample_completed_
      -- CP-element group 391: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Sample/$exit
      -- CP-element group 391: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Sample/ra
      -- 
    ra_5953_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2365_inst_ack_0, ack => convolve_CP_4675_elements(391)); -- 
    -- CP-element group 392:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 392: predecessors 
    -- CP-element group 392: 	390 
    -- CP-element group 392: successors 
    -- CP-element group 392: 	522 
    -- CP-element group 392: marked-successors 
    -- CP-element group 392: 	390 
    -- CP-element group 392: 	48 
    -- CP-element group 392: 	29 
    -- CP-element group 392:  members (3) 
      -- CP-element group 392: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_update_completed_
      -- CP-element group 392: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Update/$exit
      -- CP-element group 392: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2365_Update/ca
      -- 
    ca_5958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 392_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2365_inst_ack_1, ack => convolve_CP_4675_elements(392)); -- 
    -- CP-element group 393:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 393: predecessors 
    -- CP-element group 393: 	348 
    -- CP-element group 393: 	360 
    -- CP-element group 393: 	372 
    -- CP-element group 393: marked-predecessors 
    -- CP-element group 393: 	395 
    -- CP-element group 393: successors 
    -- CP-element group 393: 	395 
    -- CP-element group 393:  members (3) 
      -- CP-element group 393: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_sample_start_
      -- CP-element group 393: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Sample/$entry
      -- CP-element group 393: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Sample/rr
      -- 
    rr_5966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(393), ack => slice_2369_inst_req_0); -- 
    convolve_cp_element_group_393: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_393"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(395);
      gj_convolve_cp_element_group_393 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(393), clk => clk, reset => reset); --
    end block;
    -- CP-element group 394:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 394: predecessors 
    -- CP-element group 394: 	26 
    -- CP-element group 394: marked-predecessors 
    -- CP-element group 394: 	396 
    -- CP-element group 394: 	524 
    -- CP-element group 394: successors 
    -- CP-element group 394: 	396 
    -- CP-element group 394:  members (3) 
      -- CP-element group 394: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_update_start_
      -- CP-element group 394: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Update/$entry
      -- CP-element group 394: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Update/cr
      -- 
    cr_5971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(394), ack => slice_2369_inst_req_1); -- 
    convolve_cp_element_group_394: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_394"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(396) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_394 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(394), clk => clk, reset => reset); --
    end block;
    -- CP-element group 395:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 395: predecessors 
    -- CP-element group 395: 	393 
    -- CP-element group 395: successors 
    -- CP-element group 395: marked-successors 
    -- CP-element group 395: 	346 
    -- CP-element group 395: 	358 
    -- CP-element group 395: 	393 
    -- CP-element group 395: 	370 
    -- CP-element group 395:  members (3) 
      -- CP-element group 395: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_sample_completed_
      -- CP-element group 395: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Sample/$exit
      -- CP-element group 395: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Sample/ra
      -- 
    ra_5967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 395_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2369_inst_ack_0, ack => convolve_CP_4675_elements(395)); -- 
    -- CP-element group 396:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 396: predecessors 
    -- CP-element group 396: 	394 
    -- CP-element group 396: successors 
    -- CP-element group 396: 	522 
    -- CP-element group 396: marked-successors 
    -- CP-element group 396: 	48 
    -- CP-element group 396: 	394 
    -- CP-element group 396: 	29 
    -- CP-element group 396:  members (3) 
      -- CP-element group 396: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_update_completed_
      -- CP-element group 396: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Update/$exit
      -- CP-element group 396: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2369_Update/ca
      -- 
    ca_5972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 396_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2369_inst_ack_1, ack => convolve_CP_4675_elements(396)); -- 
    -- CP-element group 397:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 397: predecessors 
    -- CP-element group 397: 	348 
    -- CP-element group 397: 	360 
    -- CP-element group 397: 	372 
    -- CP-element group 397: marked-predecessors 
    -- CP-element group 397: 	399 
    -- CP-element group 397: successors 
    -- CP-element group 397: 	399 
    -- CP-element group 397:  members (3) 
      -- CP-element group 397: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_sample_start_
      -- CP-element group 397: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Sample/$entry
      -- CP-element group 397: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Sample/rr
      -- 
    rr_5980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(397), ack => slice_2373_inst_req_0); -- 
    convolve_cp_element_group_397: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_397"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(399);
      gj_convolve_cp_element_group_397 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(397), clk => clk, reset => reset); --
    end block;
    -- CP-element group 398:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 398: predecessors 
    -- CP-element group 398: 	26 
    -- CP-element group 398: marked-predecessors 
    -- CP-element group 398: 	400 
    -- CP-element group 398: 	524 
    -- CP-element group 398: successors 
    -- CP-element group 398: 	400 
    -- CP-element group 398:  members (3) 
      -- CP-element group 398: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_update_start_
      -- CP-element group 398: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Update/$entry
      -- CP-element group 398: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Update/cr
      -- 
    cr_5985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(398), ack => slice_2373_inst_req_1); -- 
    convolve_cp_element_group_398: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_398"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(400) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_398 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(398), clk => clk, reset => reset); --
    end block;
    -- CP-element group 399:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 399: predecessors 
    -- CP-element group 399: 	397 
    -- CP-element group 399: successors 
    -- CP-element group 399: marked-successors 
    -- CP-element group 399: 	346 
    -- CP-element group 399: 	358 
    -- CP-element group 399: 	370 
    -- CP-element group 399: 	397 
    -- CP-element group 399:  members (3) 
      -- CP-element group 399: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_sample_completed_
      -- CP-element group 399: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Sample/$exit
      -- CP-element group 399: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Sample/ra
      -- 
    ra_5981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 399_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2373_inst_ack_0, ack => convolve_CP_4675_elements(399)); -- 
    -- CP-element group 400:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 400: predecessors 
    -- CP-element group 400: 	398 
    -- CP-element group 400: successors 
    -- CP-element group 400: 	522 
    -- CP-element group 400: marked-successors 
    -- CP-element group 400: 	48 
    -- CP-element group 400: 	398 
    -- CP-element group 400: 	29 
    -- CP-element group 400:  members (3) 
      -- CP-element group 400: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_update_completed_
      -- CP-element group 400: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Update/$exit
      -- CP-element group 400: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2373_Update/ca
      -- 
    ca_5986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 400_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2373_inst_ack_1, ack => convolve_CP_4675_elements(400)); -- 
    -- CP-element group 401:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 401: predecessors 
    -- CP-element group 401: 	348 
    -- CP-element group 401: 	360 
    -- CP-element group 401: 	372 
    -- CP-element group 401: marked-predecessors 
    -- CP-element group 401: 	403 
    -- CP-element group 401: successors 
    -- CP-element group 401: 	403 
    -- CP-element group 401:  members (3) 
      -- CP-element group 401: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_sample_start_
      -- CP-element group 401: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Sample/$entry
      -- CP-element group 401: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Sample/rr
      -- 
    rr_5994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(401), ack => slice_2377_inst_req_0); -- 
    convolve_cp_element_group_401: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_401"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(403);
      gj_convolve_cp_element_group_401 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(401), clk => clk, reset => reset); --
    end block;
    -- CP-element group 402:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 402: predecessors 
    -- CP-element group 402: 	26 
    -- CP-element group 402: marked-predecessors 
    -- CP-element group 402: 	404 
    -- CP-element group 402: 	524 
    -- CP-element group 402: successors 
    -- CP-element group 402: 	404 
    -- CP-element group 402:  members (3) 
      -- CP-element group 402: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_update_start_
      -- CP-element group 402: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Update/$entry
      -- CP-element group 402: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Update/cr
      -- 
    cr_5999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(402), ack => slice_2377_inst_req_1); -- 
    convolve_cp_element_group_402: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_402"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(404) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_402 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(402), clk => clk, reset => reset); --
    end block;
    -- CP-element group 403:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 403: predecessors 
    -- CP-element group 403: 	401 
    -- CP-element group 403: successors 
    -- CP-element group 403: marked-successors 
    -- CP-element group 403: 	346 
    -- CP-element group 403: 	358 
    -- CP-element group 403: 	370 
    -- CP-element group 403: 	401 
    -- CP-element group 403:  members (3) 
      -- CP-element group 403: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_sample_completed_
      -- CP-element group 403: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Sample/$exit
      -- CP-element group 403: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Sample/ra
      -- 
    ra_5995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 403_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2377_inst_ack_0, ack => convolve_CP_4675_elements(403)); -- 
    -- CP-element group 404:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 404: predecessors 
    -- CP-element group 404: 	402 
    -- CP-element group 404: successors 
    -- CP-element group 404: 	522 
    -- CP-element group 404: marked-successors 
    -- CP-element group 404: 	48 
    -- CP-element group 404: 	402 
    -- CP-element group 404: 	29 
    -- CP-element group 404:  members (3) 
      -- CP-element group 404: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_update_completed_
      -- CP-element group 404: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Update/$exit
      -- CP-element group 404: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2377_Update/ca
      -- 
    ca_6000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 404_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2377_inst_ack_1, ack => convolve_CP_4675_elements(404)); -- 
    -- CP-element group 405:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 405: predecessors 
    -- CP-element group 405: 	348 
    -- CP-element group 405: 	360 
    -- CP-element group 405: 	372 
    -- CP-element group 405: marked-predecessors 
    -- CP-element group 405: 	407 
    -- CP-element group 405: successors 
    -- CP-element group 405: 	407 
    -- CP-element group 405:  members (3) 
      -- CP-element group 405: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_sample_start_
      -- CP-element group 405: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Sample/$entry
      -- CP-element group 405: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Sample/rr
      -- 
    rr_6008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(405), ack => slice_2381_inst_req_0); -- 
    convolve_cp_element_group_405: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_405"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(407);
      gj_convolve_cp_element_group_405 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(405), clk => clk, reset => reset); --
    end block;
    -- CP-element group 406:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 406: predecessors 
    -- CP-element group 406: 	26 
    -- CP-element group 406: marked-predecessors 
    -- CP-element group 406: 	408 
    -- CP-element group 406: 	524 
    -- CP-element group 406: successors 
    -- CP-element group 406: 	408 
    -- CP-element group 406:  members (3) 
      -- CP-element group 406: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_update_start_
      -- CP-element group 406: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Update/$entry
      -- CP-element group 406: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Update/cr
      -- 
    cr_6013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(406), ack => slice_2381_inst_req_1); -- 
    convolve_cp_element_group_406: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_406"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(408) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_406 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(406), clk => clk, reset => reset); --
    end block;
    -- CP-element group 407:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 407: predecessors 
    -- CP-element group 407: 	405 
    -- CP-element group 407: successors 
    -- CP-element group 407: marked-successors 
    -- CP-element group 407: 	346 
    -- CP-element group 407: 	358 
    -- CP-element group 407: 	370 
    -- CP-element group 407: 	405 
    -- CP-element group 407:  members (3) 
      -- CP-element group 407: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_sample_completed_
      -- CP-element group 407: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Sample/$exit
      -- CP-element group 407: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Sample/ra
      -- 
    ra_6009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 407_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2381_inst_ack_0, ack => convolve_CP_4675_elements(407)); -- 
    -- CP-element group 408:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 408: predecessors 
    -- CP-element group 408: 	406 
    -- CP-element group 408: successors 
    -- CP-element group 408: 	522 
    -- CP-element group 408: marked-successors 
    -- CP-element group 408: 	48 
    -- CP-element group 408: 	406 
    -- CP-element group 408: 	29 
    -- CP-element group 408:  members (3) 
      -- CP-element group 408: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_update_completed_
      -- CP-element group 408: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Update/$exit
      -- CP-element group 408: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2381_Update/ca
      -- 
    ca_6014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 408_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2381_inst_ack_1, ack => convolve_CP_4675_elements(408)); -- 
    -- CP-element group 409:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 409: predecessors 
    -- CP-element group 409: 	348 
    -- CP-element group 409: 	360 
    -- CP-element group 409: 	372 
    -- CP-element group 409: marked-predecessors 
    -- CP-element group 409: 	411 
    -- CP-element group 409: successors 
    -- CP-element group 409: 	411 
    -- CP-element group 409:  members (3) 
      -- CP-element group 409: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_sample_start_
      -- CP-element group 409: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Sample/$entry
      -- CP-element group 409: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Sample/rr
      -- 
    rr_6022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(409), ack => slice_2385_inst_req_0); -- 
    convolve_cp_element_group_409: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_409"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(411);
      gj_convolve_cp_element_group_409 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(409), clk => clk, reset => reset); --
    end block;
    -- CP-element group 410:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 410: predecessors 
    -- CP-element group 410: 	26 
    -- CP-element group 410: marked-predecessors 
    -- CP-element group 410: 	524 
    -- CP-element group 410: 	412 
    -- CP-element group 410: successors 
    -- CP-element group 410: 	412 
    -- CP-element group 410:  members (3) 
      -- CP-element group 410: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_update_start_
      -- CP-element group 410: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Update/$entry
      -- CP-element group 410: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Update/cr
      -- 
    cr_6027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(410), ack => slice_2385_inst_req_1); -- 
    convolve_cp_element_group_410: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_410"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(412);
      gj_convolve_cp_element_group_410 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(410), clk => clk, reset => reset); --
    end block;
    -- CP-element group 411:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 411: predecessors 
    -- CP-element group 411: 	409 
    -- CP-element group 411: successors 
    -- CP-element group 411: marked-successors 
    -- CP-element group 411: 	346 
    -- CP-element group 411: 	409 
    -- CP-element group 411: 	358 
    -- CP-element group 411: 	370 
    -- CP-element group 411:  members (3) 
      -- CP-element group 411: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_sample_completed_
      -- CP-element group 411: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Sample/$exit
      -- CP-element group 411: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Sample/ra
      -- 
    ra_6023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 411_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2385_inst_ack_0, ack => convolve_CP_4675_elements(411)); -- 
    -- CP-element group 412:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 412: predecessors 
    -- CP-element group 412: 	410 
    -- CP-element group 412: successors 
    -- CP-element group 412: 	522 
    -- CP-element group 412: marked-successors 
    -- CP-element group 412: 	410 
    -- CP-element group 412: 	48 
    -- CP-element group 412: 	29 
    -- CP-element group 412:  members (3) 
      -- CP-element group 412: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_update_completed_
      -- CP-element group 412: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Update/$exit
      -- CP-element group 412: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2385_Update/ca
      -- 
    ca_6028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 412_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2385_inst_ack_1, ack => convolve_CP_4675_elements(412)); -- 
    -- CP-element group 413:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 413: predecessors 
    -- CP-element group 413: 	352 
    -- CP-element group 413: 	364 
    -- CP-element group 413: 	376 
    -- CP-element group 413: marked-predecessors 
    -- CP-element group 413: 	415 
    -- CP-element group 413: successors 
    -- CP-element group 413: 	415 
    -- CP-element group 413:  members (3) 
      -- CP-element group 413: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_sample_start_
      -- CP-element group 413: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Sample/$entry
      -- CP-element group 413: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Sample/rr
      -- 
    rr_6036_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6036_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(413), ack => slice_2389_inst_req_0); -- 
    convolve_cp_element_group_413: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_413"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(415);
      gj_convolve_cp_element_group_413 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(413), clk => clk, reset => reset); --
    end block;
    -- CP-element group 414:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 414: predecessors 
    -- CP-element group 414: 	26 
    -- CP-element group 414: marked-predecessors 
    -- CP-element group 414: 	524 
    -- CP-element group 414: 	416 
    -- CP-element group 414: successors 
    -- CP-element group 414: 	416 
    -- CP-element group 414:  members (3) 
      -- CP-element group 414: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_update_start_
      -- CP-element group 414: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Update/$entry
      -- CP-element group 414: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Update/cr
      -- 
    cr_6041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(414), ack => slice_2389_inst_req_1); -- 
    convolve_cp_element_group_414: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_414"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(416);
      gj_convolve_cp_element_group_414 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(414), clk => clk, reset => reset); --
    end block;
    -- CP-element group 415:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 415: predecessors 
    -- CP-element group 415: 	413 
    -- CP-element group 415: successors 
    -- CP-element group 415: marked-successors 
    -- CP-element group 415: 	362 
    -- CP-element group 415: 	350 
    -- CP-element group 415: 	374 
    -- CP-element group 415: 	413 
    -- CP-element group 415:  members (3) 
      -- CP-element group 415: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_sample_completed_
      -- CP-element group 415: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Sample/$exit
      -- CP-element group 415: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Sample/ra
      -- 
    ra_6037_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 415_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2389_inst_ack_0, ack => convolve_CP_4675_elements(415)); -- 
    -- CP-element group 416:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 416: predecessors 
    -- CP-element group 416: 	414 
    -- CP-element group 416: successors 
    -- CP-element group 416: 	522 
    -- CP-element group 416: marked-successors 
    -- CP-element group 416: 	48 
    -- CP-element group 416: 	29 
    -- CP-element group 416: 	414 
    -- CP-element group 416:  members (3) 
      -- CP-element group 416: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_update_completed_
      -- CP-element group 416: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Update/$exit
      -- CP-element group 416: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2389_Update/ca
      -- 
    ca_6042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 416_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2389_inst_ack_1, ack => convolve_CP_4675_elements(416)); -- 
    -- CP-element group 417:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 417: predecessors 
    -- CP-element group 417: 	352 
    -- CP-element group 417: 	364 
    -- CP-element group 417: 	376 
    -- CP-element group 417: marked-predecessors 
    -- CP-element group 417: 	419 
    -- CP-element group 417: successors 
    -- CP-element group 417: 	419 
    -- CP-element group 417:  members (3) 
      -- CP-element group 417: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_sample_start_
      -- CP-element group 417: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Sample/$entry
      -- CP-element group 417: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Sample/rr
      -- 
    rr_6050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(417), ack => slice_2393_inst_req_0); -- 
    convolve_cp_element_group_417: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_417"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(419);
      gj_convolve_cp_element_group_417 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(417), clk => clk, reset => reset); --
    end block;
    -- CP-element group 418:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 418: predecessors 
    -- CP-element group 418: 	26 
    -- CP-element group 418: marked-predecessors 
    -- CP-element group 418: 	420 
    -- CP-element group 418: 	524 
    -- CP-element group 418: successors 
    -- CP-element group 418: 	420 
    -- CP-element group 418:  members (3) 
      -- CP-element group 418: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_update_start_
      -- CP-element group 418: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Update/$entry
      -- CP-element group 418: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Update/cr
      -- 
    cr_6055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(418), ack => slice_2393_inst_req_1); -- 
    convolve_cp_element_group_418: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_418"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(420) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_418 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(418), clk => clk, reset => reset); --
    end block;
    -- CP-element group 419:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 419: predecessors 
    -- CP-element group 419: 	417 
    -- CP-element group 419: successors 
    -- CP-element group 419: marked-successors 
    -- CP-element group 419: 	362 
    -- CP-element group 419: 	350 
    -- CP-element group 419: 	374 
    -- CP-element group 419: 	417 
    -- CP-element group 419:  members (3) 
      -- CP-element group 419: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_sample_completed_
      -- CP-element group 419: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Sample/$exit
      -- CP-element group 419: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Sample/ra
      -- 
    ra_6051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 419_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2393_inst_ack_0, ack => convolve_CP_4675_elements(419)); -- 
    -- CP-element group 420:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 420: predecessors 
    -- CP-element group 420: 	418 
    -- CP-element group 420: successors 
    -- CP-element group 420: 	522 
    -- CP-element group 420: marked-successors 
    -- CP-element group 420: 	48 
    -- CP-element group 420: 	29 
    -- CP-element group 420: 	418 
    -- CP-element group 420:  members (3) 
      -- CP-element group 420: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_update_completed_
      -- CP-element group 420: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Update/$exit
      -- CP-element group 420: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2393_Update/ca
      -- 
    ca_6056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 420_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2393_inst_ack_1, ack => convolve_CP_4675_elements(420)); -- 
    -- CP-element group 421:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 421: predecessors 
    -- CP-element group 421: 	352 
    -- CP-element group 421: 	364 
    -- CP-element group 421: 	376 
    -- CP-element group 421: marked-predecessors 
    -- CP-element group 421: 	423 
    -- CP-element group 421: successors 
    -- CP-element group 421: 	423 
    -- CP-element group 421:  members (3) 
      -- CP-element group 421: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Sample/rr
      -- CP-element group 421: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Sample/$entry
      -- CP-element group 421: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_sample_start_
      -- 
    rr_6064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(421), ack => slice_2397_inst_req_0); -- 
    convolve_cp_element_group_421: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_421"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(423);
      gj_convolve_cp_element_group_421 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(421), clk => clk, reset => reset); --
    end block;
    -- CP-element group 422:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 422: predecessors 
    -- CP-element group 422: 	26 
    -- CP-element group 422: marked-predecessors 
    -- CP-element group 422: 	424 
    -- CP-element group 422: 	524 
    -- CP-element group 422: successors 
    -- CP-element group 422: 	424 
    -- CP-element group 422:  members (3) 
      -- CP-element group 422: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Update/cr
      -- CP-element group 422: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Update/$entry
      -- CP-element group 422: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_update_start_
      -- 
    cr_6069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(422), ack => slice_2397_inst_req_1); -- 
    convolve_cp_element_group_422: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_422"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(424) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_422 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(422), clk => clk, reset => reset); --
    end block;
    -- CP-element group 423:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 423: predecessors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: successors 
    -- CP-element group 423: marked-successors 
    -- CP-element group 423: 	421 
    -- CP-element group 423: 	362 
    -- CP-element group 423: 	350 
    -- CP-element group 423: 	374 
    -- CP-element group 423:  members (3) 
      -- CP-element group 423: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Sample/ra
      -- CP-element group 423: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Sample/$exit
      -- CP-element group 423: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_sample_completed_
      -- 
    ra_6065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 423_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2397_inst_ack_0, ack => convolve_CP_4675_elements(423)); -- 
    -- CP-element group 424:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 424: predecessors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: successors 
    -- CP-element group 424: 	522 
    -- CP-element group 424: marked-successors 
    -- CP-element group 424: 	422 
    -- CP-element group 424: 	48 
    -- CP-element group 424: 	29 
    -- CP-element group 424:  members (3) 
      -- CP-element group 424: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Update/ca
      -- CP-element group 424: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_Update/$exit
      -- CP-element group 424: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2397_update_completed_
      -- 
    ca_6070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 424_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2397_inst_ack_1, ack => convolve_CP_4675_elements(424)); -- 
    -- CP-element group 425:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 425: predecessors 
    -- CP-element group 425: 	352 
    -- CP-element group 425: 	364 
    -- CP-element group 425: 	376 
    -- CP-element group 425: marked-predecessors 
    -- CP-element group 425: 	427 
    -- CP-element group 425: successors 
    -- CP-element group 425: 	427 
    -- CP-element group 425:  members (3) 
      -- CP-element group 425: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_sample_start_
      -- CP-element group 425: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Sample/$entry
      -- CP-element group 425: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Sample/rr
      -- 
    rr_6078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(425), ack => slice_2401_inst_req_0); -- 
    convolve_cp_element_group_425: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_425"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(427);
      gj_convolve_cp_element_group_425 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(425), clk => clk, reset => reset); --
    end block;
    -- CP-element group 426:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 426: predecessors 
    -- CP-element group 426: 	26 
    -- CP-element group 426: marked-predecessors 
    -- CP-element group 426: 	428 
    -- CP-element group 426: 	524 
    -- CP-element group 426: successors 
    -- CP-element group 426: 	428 
    -- CP-element group 426:  members (3) 
      -- CP-element group 426: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_update_start_
      -- CP-element group 426: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Update/$entry
      -- CP-element group 426: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Update/cr
      -- 
    cr_6083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(426), ack => slice_2401_inst_req_1); -- 
    convolve_cp_element_group_426: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_426"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(428) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_426 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(426), clk => clk, reset => reset); --
    end block;
    -- CP-element group 427:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 427: predecessors 
    -- CP-element group 427: 	425 
    -- CP-element group 427: successors 
    -- CP-element group 427: marked-successors 
    -- CP-element group 427: 	362 
    -- CP-element group 427: 	350 
    -- CP-element group 427: 	374 
    -- CP-element group 427: 	425 
    -- CP-element group 427:  members (3) 
      -- CP-element group 427: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_sample_completed_
      -- CP-element group 427: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Sample/$exit
      -- CP-element group 427: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Sample/ra
      -- 
    ra_6079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 427_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2401_inst_ack_0, ack => convolve_CP_4675_elements(427)); -- 
    -- CP-element group 428:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 428: predecessors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: successors 
    -- CP-element group 428: 	522 
    -- CP-element group 428: marked-successors 
    -- CP-element group 428: 	426 
    -- CP-element group 428: 	48 
    -- CP-element group 428: 	29 
    -- CP-element group 428:  members (3) 
      -- CP-element group 428: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_update_completed_
      -- CP-element group 428: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Update/$exit
      -- CP-element group 428: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2401_Update/ca
      -- 
    ca_6084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 428_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2401_inst_ack_1, ack => convolve_CP_4675_elements(428)); -- 
    -- CP-element group 429:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 429: predecessors 
    -- CP-element group 429: 	352 
    -- CP-element group 429: 	364 
    -- CP-element group 429: 	376 
    -- CP-element group 429: marked-predecessors 
    -- CP-element group 429: 	431 
    -- CP-element group 429: successors 
    -- CP-element group 429: 	431 
    -- CP-element group 429:  members (3) 
      -- CP-element group 429: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Sample/$entry
      -- CP-element group 429: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Sample/rr
      -- CP-element group 429: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_sample_start_
      -- 
    rr_6092_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6092_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(429), ack => slice_2405_inst_req_0); -- 
    convolve_cp_element_group_429: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_429"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(431);
      gj_convolve_cp_element_group_429 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(429), clk => clk, reset => reset); --
    end block;
    -- CP-element group 430:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 430: predecessors 
    -- CP-element group 430: 	26 
    -- CP-element group 430: marked-predecessors 
    -- CP-element group 430: 	524 
    -- CP-element group 430: 	432 
    -- CP-element group 430: successors 
    -- CP-element group 430: 	432 
    -- CP-element group 430:  members (3) 
      -- CP-element group 430: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_update_start_
      -- CP-element group 430: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Update/$entry
      -- CP-element group 430: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Update/cr
      -- 
    cr_6097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(430), ack => slice_2405_inst_req_1); -- 
    convolve_cp_element_group_430: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_430"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(432);
      gj_convolve_cp_element_group_430 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(430), clk => clk, reset => reset); --
    end block;
    -- CP-element group 431:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 431: predecessors 
    -- CP-element group 431: 	429 
    -- CP-element group 431: successors 
    -- CP-element group 431: marked-successors 
    -- CP-element group 431: 	362 
    -- CP-element group 431: 	350 
    -- CP-element group 431: 	374 
    -- CP-element group 431: 	429 
    -- CP-element group 431:  members (3) 
      -- CP-element group 431: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_sample_completed_
      -- CP-element group 431: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Sample/$exit
      -- CP-element group 431: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Sample/ra
      -- 
    ra_6093_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 431_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2405_inst_ack_0, ack => convolve_CP_4675_elements(431)); -- 
    -- CP-element group 432:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 432: predecessors 
    -- CP-element group 432: 	430 
    -- CP-element group 432: successors 
    -- CP-element group 432: 	522 
    -- CP-element group 432: marked-successors 
    -- CP-element group 432: 	430 
    -- CP-element group 432: 	48 
    -- CP-element group 432: 	29 
    -- CP-element group 432:  members (3) 
      -- CP-element group 432: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_update_completed_
      -- CP-element group 432: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Update/$exit
      -- CP-element group 432: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2405_Update/ca
      -- 
    ca_6098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 432_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2405_inst_ack_1, ack => convolve_CP_4675_elements(432)); -- 
    -- CP-element group 433:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 433: predecessors 
    -- CP-element group 433: 	352 
    -- CP-element group 433: 	364 
    -- CP-element group 433: 	376 
    -- CP-element group 433: marked-predecessors 
    -- CP-element group 433: 	435 
    -- CP-element group 433: successors 
    -- CP-element group 433: 	435 
    -- CP-element group 433:  members (3) 
      -- CP-element group 433: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Sample/rr
      -- CP-element group 433: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Sample/$entry
      -- CP-element group 433: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_sample_start_
      -- 
    rr_6106_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6106_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(433), ack => slice_2409_inst_req_0); -- 
    convolve_cp_element_group_433: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_433"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(435);
      gj_convolve_cp_element_group_433 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(433), clk => clk, reset => reset); --
    end block;
    -- CP-element group 434:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 434: predecessors 
    -- CP-element group 434: 	26 
    -- CP-element group 434: marked-predecessors 
    -- CP-element group 434: 	436 
    -- CP-element group 434: 	524 
    -- CP-element group 434: successors 
    -- CP-element group 434: 	436 
    -- CP-element group 434:  members (3) 
      -- CP-element group 434: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Update/cr
      -- CP-element group 434: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Update/$entry
      -- CP-element group 434: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_update_start_
      -- 
    cr_6111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(434), ack => slice_2409_inst_req_1); -- 
    convolve_cp_element_group_434: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_434"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(436) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_434 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(434), clk => clk, reset => reset); --
    end block;
    -- CP-element group 435:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 435: predecessors 
    -- CP-element group 435: 	433 
    -- CP-element group 435: successors 
    -- CP-element group 435: marked-successors 
    -- CP-element group 435: 	362 
    -- CP-element group 435: 	350 
    -- CP-element group 435: 	374 
    -- CP-element group 435: 	433 
    -- CP-element group 435:  members (3) 
      -- CP-element group 435: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Sample/ra
      -- CP-element group 435: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Sample/$exit
      -- CP-element group 435: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_sample_completed_
      -- 
    ra_6107_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 435_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2409_inst_ack_0, ack => convolve_CP_4675_elements(435)); -- 
    -- CP-element group 436:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 436: predecessors 
    -- CP-element group 436: 	434 
    -- CP-element group 436: successors 
    -- CP-element group 436: 	522 
    -- CP-element group 436: marked-successors 
    -- CP-element group 436: 	48 
    -- CP-element group 436: 	29 
    -- CP-element group 436: 	434 
    -- CP-element group 436:  members (3) 
      -- CP-element group 436: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Update/ca
      -- CP-element group 436: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_Update/$exit
      -- CP-element group 436: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2409_update_completed_
      -- 
    ca_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 436_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2409_inst_ack_1, ack => convolve_CP_4675_elements(436)); -- 
    -- CP-element group 437:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 437: predecessors 
    -- CP-element group 437: 	352 
    -- CP-element group 437: 	364 
    -- CP-element group 437: 	376 
    -- CP-element group 437: marked-predecessors 
    -- CP-element group 437: 	439 
    -- CP-element group 437: successors 
    -- CP-element group 437: 	439 
    -- CP-element group 437:  members (3) 
      -- CP-element group 437: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Sample/$entry
      -- CP-element group 437: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Sample/rr
      -- CP-element group 437: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_sample_start_
      -- 
    rr_6120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(437), ack => slice_2413_inst_req_0); -- 
    convolve_cp_element_group_437: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_437"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(439);
      gj_convolve_cp_element_group_437 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(437), clk => clk, reset => reset); --
    end block;
    -- CP-element group 438:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 438: predecessors 
    -- CP-element group 438: 	26 
    -- CP-element group 438: marked-predecessors 
    -- CP-element group 438: 	440 
    -- CP-element group 438: 	524 
    -- CP-element group 438: successors 
    -- CP-element group 438: 	440 
    -- CP-element group 438:  members (3) 
      -- CP-element group 438: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_update_start_
      -- CP-element group 438: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Update/$entry
      -- CP-element group 438: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Update/cr
      -- 
    cr_6125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(438), ack => slice_2413_inst_req_1); -- 
    convolve_cp_element_group_438: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_438"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(440) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_438 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(438), clk => clk, reset => reset); --
    end block;
    -- CP-element group 439:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 439: predecessors 
    -- CP-element group 439: 	437 
    -- CP-element group 439: successors 
    -- CP-element group 439: marked-successors 
    -- CP-element group 439: 	437 
    -- CP-element group 439: 	362 
    -- CP-element group 439: 	350 
    -- CP-element group 439: 	374 
    -- CP-element group 439:  members (3) 
      -- CP-element group 439: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_sample_completed_
      -- CP-element group 439: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Sample/$exit
      -- CP-element group 439: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Sample/ra
      -- 
    ra_6121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 439_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2413_inst_ack_0, ack => convolve_CP_4675_elements(439)); -- 
    -- CP-element group 440:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 440: predecessors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: successors 
    -- CP-element group 440: 	522 
    -- CP-element group 440: marked-successors 
    -- CP-element group 440: 	438 
    -- CP-element group 440: 	48 
    -- CP-element group 440: 	29 
    -- CP-element group 440:  members (3) 
      -- CP-element group 440: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_update_completed_
      -- CP-element group 440: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Update/$exit
      -- CP-element group 440: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2413_Update/ca
      -- 
    ca_6126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 440_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2413_inst_ack_1, ack => convolve_CP_4675_elements(440)); -- 
    -- CP-element group 441:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 441: predecessors 
    -- CP-element group 441: 	352 
    -- CP-element group 441: 	364 
    -- CP-element group 441: 	376 
    -- CP-element group 441: marked-predecessors 
    -- CP-element group 441: 	443 
    -- CP-element group 441: successors 
    -- CP-element group 441: 	443 
    -- CP-element group 441:  members (3) 
      -- CP-element group 441: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_sample_start_
      -- CP-element group 441: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Sample/$entry
      -- CP-element group 441: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Sample/rr
      -- 
    rr_6134_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6134_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(441), ack => slice_2417_inst_req_0); -- 
    convolve_cp_element_group_441: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_441"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(443);
      gj_convolve_cp_element_group_441 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(441), clk => clk, reset => reset); --
    end block;
    -- CP-element group 442:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 442: predecessors 
    -- CP-element group 442: 	26 
    -- CP-element group 442: marked-predecessors 
    -- CP-element group 442: 	444 
    -- CP-element group 442: 	524 
    -- CP-element group 442: successors 
    -- CP-element group 442: 	444 
    -- CP-element group 442:  members (3) 
      -- CP-element group 442: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_update_start_
      -- CP-element group 442: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Update/$entry
      -- CP-element group 442: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Update/cr
      -- 
    cr_6139_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6139_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(442), ack => slice_2417_inst_req_1); -- 
    convolve_cp_element_group_442: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_442"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(444) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_442 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(442), clk => clk, reset => reset); --
    end block;
    -- CP-element group 443:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 443: predecessors 
    -- CP-element group 443: 	441 
    -- CP-element group 443: successors 
    -- CP-element group 443: marked-successors 
    -- CP-element group 443: 	441 
    -- CP-element group 443: 	362 
    -- CP-element group 443: 	350 
    -- CP-element group 443: 	374 
    -- CP-element group 443:  members (3) 
      -- CP-element group 443: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_sample_completed_
      -- CP-element group 443: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Sample/$exit
      -- CP-element group 443: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Sample/ra
      -- 
    ra_6135_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 443_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2417_inst_ack_0, ack => convolve_CP_4675_elements(443)); -- 
    -- CP-element group 444:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 444: predecessors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: successors 
    -- CP-element group 444: 	522 
    -- CP-element group 444: marked-successors 
    -- CP-element group 444: 	442 
    -- CP-element group 444: 	48 
    -- CP-element group 444: 	29 
    -- CP-element group 444:  members (3) 
      -- CP-element group 444: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_update_completed_
      -- CP-element group 444: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Update/$exit
      -- CP-element group 444: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2417_Update/ca
      -- 
    ca_6140_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 444_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2417_inst_ack_1, ack => convolve_CP_4675_elements(444)); -- 
    -- CP-element group 445:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 445: predecessors 
    -- CP-element group 445: 	356 
    -- CP-element group 445: 	368 
    -- CP-element group 445: 	380 
    -- CP-element group 445: marked-predecessors 
    -- CP-element group 445: 	447 
    -- CP-element group 445: successors 
    -- CP-element group 445: 	447 
    -- CP-element group 445:  members (3) 
      -- CP-element group 445: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_sample_start_
      -- CP-element group 445: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Sample/rr
      -- CP-element group 445: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Sample/$entry
      -- 
    rr_6148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(445), ack => slice_2421_inst_req_0); -- 
    convolve_cp_element_group_445: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_445"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(447);
      gj_convolve_cp_element_group_445 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(445), clk => clk, reset => reset); --
    end block;
    -- CP-element group 446:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 446: predecessors 
    -- CP-element group 446: 	26 
    -- CP-element group 446: marked-predecessors 
    -- CP-element group 446: 	448 
    -- CP-element group 446: 	524 
    -- CP-element group 446: successors 
    -- CP-element group 446: 	448 
    -- CP-element group 446:  members (3) 
      -- CP-element group 446: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_update_start_
      -- CP-element group 446: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Update/cr
      -- CP-element group 446: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Update/$entry
      -- 
    cr_6153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(446), ack => slice_2421_inst_req_1); -- 
    convolve_cp_element_group_446: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_446"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(448) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_446 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(446), clk => clk, reset => reset); --
    end block;
    -- CP-element group 447:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 447: predecessors 
    -- CP-element group 447: 	445 
    -- CP-element group 447: successors 
    -- CP-element group 447: marked-successors 
    -- CP-element group 447: 	445 
    -- CP-element group 447: 	354 
    -- CP-element group 447: 	366 
    -- CP-element group 447: 	378 
    -- CP-element group 447:  members (3) 
      -- CP-element group 447: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_sample_completed_
      -- CP-element group 447: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Sample/ra
      -- CP-element group 447: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Sample/$exit
      -- 
    ra_6149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 447_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2421_inst_ack_0, ack => convolve_CP_4675_elements(447)); -- 
    -- CP-element group 448:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 448: predecessors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: successors 
    -- CP-element group 448: 	522 
    -- CP-element group 448: marked-successors 
    -- CP-element group 448: 	446 
    -- CP-element group 448: 	48 
    -- CP-element group 448: 	29 
    -- CP-element group 448:  members (3) 
      -- CP-element group 448: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_update_completed_
      -- CP-element group 448: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Update/ca
      -- CP-element group 448: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2421_Update/$exit
      -- 
    ca_6154_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 448_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2421_inst_ack_1, ack => convolve_CP_4675_elements(448)); -- 
    -- CP-element group 449:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 449: predecessors 
    -- CP-element group 449: 	356 
    -- CP-element group 449: 	368 
    -- CP-element group 449: 	380 
    -- CP-element group 449: marked-predecessors 
    -- CP-element group 449: 	451 
    -- CP-element group 449: successors 
    -- CP-element group 449: 	451 
    -- CP-element group 449:  members (3) 
      -- CP-element group 449: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Sample/$entry
      -- CP-element group 449: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Sample/rr
      -- CP-element group 449: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_sample_start_
      -- 
    rr_6162_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6162_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(449), ack => slice_2425_inst_req_0); -- 
    convolve_cp_element_group_449: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_449"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(451);
      gj_convolve_cp_element_group_449 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(449), clk => clk, reset => reset); --
    end block;
    -- CP-element group 450:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 450: predecessors 
    -- CP-element group 450: 	26 
    -- CP-element group 450: marked-predecessors 
    -- CP-element group 450: 	452 
    -- CP-element group 450: 	524 
    -- CP-element group 450: successors 
    -- CP-element group 450: 	452 
    -- CP-element group 450:  members (3) 
      -- CP-element group 450: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Update/$entry
      -- CP-element group 450: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Update/cr
      -- CP-element group 450: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_update_start_
      -- 
    cr_6167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(450), ack => slice_2425_inst_req_1); -- 
    convolve_cp_element_group_450: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_450"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(452) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_450 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(450), clk => clk, reset => reset); --
    end block;
    -- CP-element group 451:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 451: predecessors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: successors 
    -- CP-element group 451: marked-successors 
    -- CP-element group 451: 	449 
    -- CP-element group 451: 	354 
    -- CP-element group 451: 	366 
    -- CP-element group 451: 	378 
    -- CP-element group 451:  members (3) 
      -- CP-element group 451: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Sample/$exit
      -- CP-element group 451: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Sample/ra
      -- CP-element group 451: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_sample_completed_
      -- 
    ra_6163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 451_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2425_inst_ack_0, ack => convolve_CP_4675_elements(451)); -- 
    -- CP-element group 452:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 452: predecessors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: successors 
    -- CP-element group 452: 	522 
    -- CP-element group 452: marked-successors 
    -- CP-element group 452: 	450 
    -- CP-element group 452: 	48 
    -- CP-element group 452: 	29 
    -- CP-element group 452:  members (3) 
      -- CP-element group 452: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_update_completed_
      -- CP-element group 452: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Update/$exit
      -- CP-element group 452: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2425_Update/ca
      -- 
    ca_6168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 452_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2425_inst_ack_1, ack => convolve_CP_4675_elements(452)); -- 
    -- CP-element group 453:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 453: predecessors 
    -- CP-element group 453: 	356 
    -- CP-element group 453: 	368 
    -- CP-element group 453: 	380 
    -- CP-element group 453: marked-predecessors 
    -- CP-element group 453: 	455 
    -- CP-element group 453: successors 
    -- CP-element group 453: 	455 
    -- CP-element group 453:  members (3) 
      -- CP-element group 453: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_sample_start_
      -- CP-element group 453: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Sample/$entry
      -- CP-element group 453: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Sample/rr
      -- 
    rr_6176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(453), ack => slice_2429_inst_req_0); -- 
    convolve_cp_element_group_453: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_453"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(455);
      gj_convolve_cp_element_group_453 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(453), clk => clk, reset => reset); --
    end block;
    -- CP-element group 454:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 454: predecessors 
    -- CP-element group 454: 	26 
    -- CP-element group 454: marked-predecessors 
    -- CP-element group 454: 	456 
    -- CP-element group 454: 	524 
    -- CP-element group 454: successors 
    -- CP-element group 454: 	456 
    -- CP-element group 454:  members (3) 
      -- CP-element group 454: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_update_start_
      -- CP-element group 454: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Update/$entry
      -- CP-element group 454: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Update/cr
      -- 
    cr_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(454), ack => slice_2429_inst_req_1); -- 
    convolve_cp_element_group_454: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_454"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(456) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_454 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(454), clk => clk, reset => reset); --
    end block;
    -- CP-element group 455:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 455: predecessors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: successors 
    -- CP-element group 455: marked-successors 
    -- CP-element group 455: 	453 
    -- CP-element group 455: 	354 
    -- CP-element group 455: 	366 
    -- CP-element group 455: 	378 
    -- CP-element group 455:  members (3) 
      -- CP-element group 455: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_sample_completed_
      -- CP-element group 455: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Sample/$exit
      -- CP-element group 455: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Sample/ra
      -- 
    ra_6177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 455_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2429_inst_ack_0, ack => convolve_CP_4675_elements(455)); -- 
    -- CP-element group 456:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 456: predecessors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: successors 
    -- CP-element group 456: 	522 
    -- CP-element group 456: marked-successors 
    -- CP-element group 456: 	454 
    -- CP-element group 456: 	48 
    -- CP-element group 456: 	29 
    -- CP-element group 456:  members (3) 
      -- CP-element group 456: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_update_completed_
      -- CP-element group 456: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Update/$exit
      -- CP-element group 456: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2429_Update/ca
      -- 
    ca_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 456_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2429_inst_ack_1, ack => convolve_CP_4675_elements(456)); -- 
    -- CP-element group 457:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 457: predecessors 
    -- CP-element group 457: 	356 
    -- CP-element group 457: 	368 
    -- CP-element group 457: 	380 
    -- CP-element group 457: marked-predecessors 
    -- CP-element group 457: 	459 
    -- CP-element group 457: successors 
    -- CP-element group 457: 	459 
    -- CP-element group 457:  members (3) 
      -- CP-element group 457: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_sample_start_
      -- CP-element group 457: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Sample/$entry
      -- CP-element group 457: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Sample/rr
      -- 
    rr_6190_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6190_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(457), ack => slice_2433_inst_req_0); -- 
    convolve_cp_element_group_457: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_457"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(459);
      gj_convolve_cp_element_group_457 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(457), clk => clk, reset => reset); --
    end block;
    -- CP-element group 458:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 458: predecessors 
    -- CP-element group 458: 	26 
    -- CP-element group 458: marked-predecessors 
    -- CP-element group 458: 	460 
    -- CP-element group 458: 	524 
    -- CP-element group 458: successors 
    -- CP-element group 458: 	460 
    -- CP-element group 458:  members (3) 
      -- CP-element group 458: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_update_start_
      -- CP-element group 458: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Update/cr
      -- CP-element group 458: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Update/$entry
      -- 
    cr_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(458), ack => slice_2433_inst_req_1); -- 
    convolve_cp_element_group_458: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_458"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(460) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_458 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(458), clk => clk, reset => reset); --
    end block;
    -- CP-element group 459:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 459: predecessors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: successors 
    -- CP-element group 459: marked-successors 
    -- CP-element group 459: 	457 
    -- CP-element group 459: 	354 
    -- CP-element group 459: 	366 
    -- CP-element group 459: 	378 
    -- CP-element group 459:  members (3) 
      -- CP-element group 459: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_sample_completed_
      -- CP-element group 459: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Sample/ra
      -- CP-element group 459: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Sample/$exit
      -- 
    ra_6191_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 459_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2433_inst_ack_0, ack => convolve_CP_4675_elements(459)); -- 
    -- CP-element group 460:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 460: predecessors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: successors 
    -- CP-element group 460: 	522 
    -- CP-element group 460: marked-successors 
    -- CP-element group 460: 	458 
    -- CP-element group 460: 	48 
    -- CP-element group 460: 	29 
    -- CP-element group 460:  members (3) 
      -- CP-element group 460: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_update_completed_
      -- CP-element group 460: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Update/ca
      -- CP-element group 460: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2433_Update/$exit
      -- 
    ca_6196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 460_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2433_inst_ack_1, ack => convolve_CP_4675_elements(460)); -- 
    -- CP-element group 461:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 461: predecessors 
    -- CP-element group 461: 	356 
    -- CP-element group 461: 	368 
    -- CP-element group 461: 	380 
    -- CP-element group 461: marked-predecessors 
    -- CP-element group 461: 	463 
    -- CP-element group 461: successors 
    -- CP-element group 461: 	463 
    -- CP-element group 461:  members (3) 
      -- CP-element group 461: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Sample/rr
      -- CP-element group 461: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Sample/$entry
      -- CP-element group 461: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_sample_start_
      -- 
    rr_6204_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6204_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(461), ack => slice_2437_inst_req_0); -- 
    convolve_cp_element_group_461: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_461"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(463);
      gj_convolve_cp_element_group_461 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(461), clk => clk, reset => reset); --
    end block;
    -- CP-element group 462:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 462: predecessors 
    -- CP-element group 462: 	26 
    -- CP-element group 462: marked-predecessors 
    -- CP-element group 462: 	464 
    -- CP-element group 462: 	524 
    -- CP-element group 462: successors 
    -- CP-element group 462: 	464 
    -- CP-element group 462:  members (3) 
      -- CP-element group 462: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Update/$entry
      -- CP-element group 462: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Update/cr
      -- CP-element group 462: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_update_start_
      -- 
    cr_6209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(462), ack => slice_2437_inst_req_1); -- 
    convolve_cp_element_group_462: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_462"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(464) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_462 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(462), clk => clk, reset => reset); --
    end block;
    -- CP-element group 463:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 463: predecessors 
    -- CP-element group 463: 	461 
    -- CP-element group 463: successors 
    -- CP-element group 463: marked-successors 
    -- CP-element group 463: 	461 
    -- CP-element group 463: 	354 
    -- CP-element group 463: 	366 
    -- CP-element group 463: 	378 
    -- CP-element group 463:  members (3) 
      -- CP-element group 463: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Sample/ra
      -- CP-element group 463: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Sample/$exit
      -- CP-element group 463: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_sample_completed_
      -- 
    ra_6205_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 463_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2437_inst_ack_0, ack => convolve_CP_4675_elements(463)); -- 
    -- CP-element group 464:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 464: predecessors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: successors 
    -- CP-element group 464: 	522 
    -- CP-element group 464: marked-successors 
    -- CP-element group 464: 	462 
    -- CP-element group 464: 	48 
    -- CP-element group 464: 	29 
    -- CP-element group 464:  members (3) 
      -- CP-element group 464: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Update/$exit
      -- CP-element group 464: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_Update/ca
      -- CP-element group 464: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2437_update_completed_
      -- 
    ca_6210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 464_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2437_inst_ack_1, ack => convolve_CP_4675_elements(464)); -- 
    -- CP-element group 465:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 465: predecessors 
    -- CP-element group 465: 	356 
    -- CP-element group 465: 	368 
    -- CP-element group 465: 	380 
    -- CP-element group 465: marked-predecessors 
    -- CP-element group 465: 	467 
    -- CP-element group 465: successors 
    -- CP-element group 465: 	467 
    -- CP-element group 465:  members (3) 
      -- CP-element group 465: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_sample_start_
      -- CP-element group 465: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Sample/$entry
      -- CP-element group 465: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Sample/rr
      -- 
    rr_6218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(465), ack => slice_2441_inst_req_0); -- 
    convolve_cp_element_group_465: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_465"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(467);
      gj_convolve_cp_element_group_465 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(465), clk => clk, reset => reset); --
    end block;
    -- CP-element group 466:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 466: predecessors 
    -- CP-element group 466: 	26 
    -- CP-element group 466: marked-predecessors 
    -- CP-element group 466: 	468 
    -- CP-element group 466: 	524 
    -- CP-element group 466: successors 
    -- CP-element group 466: 	468 
    -- CP-element group 466:  members (3) 
      -- CP-element group 466: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_update_start_
      -- CP-element group 466: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Update/$entry
      -- CP-element group 466: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Update/cr
      -- 
    cr_6223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(466), ack => slice_2441_inst_req_1); -- 
    convolve_cp_element_group_466: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_466"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(468) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_466 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(466), clk => clk, reset => reset); --
    end block;
    -- CP-element group 467:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 467: predecessors 
    -- CP-element group 467: 	465 
    -- CP-element group 467: successors 
    -- CP-element group 467: marked-successors 
    -- CP-element group 467: 	465 
    -- CP-element group 467: 	354 
    -- CP-element group 467: 	366 
    -- CP-element group 467: 	378 
    -- CP-element group 467:  members (3) 
      -- CP-element group 467: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_sample_completed_
      -- CP-element group 467: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Sample/$exit
      -- CP-element group 467: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Sample/ra
      -- 
    ra_6219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 467_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2441_inst_ack_0, ack => convolve_CP_4675_elements(467)); -- 
    -- CP-element group 468:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 468: predecessors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: successors 
    -- CP-element group 468: 	522 
    -- CP-element group 468: marked-successors 
    -- CP-element group 468: 	466 
    -- CP-element group 468: 	48 
    -- CP-element group 468: 	29 
    -- CP-element group 468:  members (3) 
      -- CP-element group 468: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_update_completed_
      -- CP-element group 468: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Update/$exit
      -- CP-element group 468: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2441_Update/ca
      -- 
    ca_6224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 468_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2441_inst_ack_1, ack => convolve_CP_4675_elements(468)); -- 
    -- CP-element group 469:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 469: predecessors 
    -- CP-element group 469: 	356 
    -- CP-element group 469: 	368 
    -- CP-element group 469: 	380 
    -- CP-element group 469: marked-predecessors 
    -- CP-element group 469: 	471 
    -- CP-element group 469: successors 
    -- CP-element group 469: 	471 
    -- CP-element group 469:  members (3) 
      -- CP-element group 469: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Sample/rr
      -- CP-element group 469: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_sample_start_
      -- CP-element group 469: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Sample/$entry
      -- 
    rr_6232_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6232_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(469), ack => slice_2445_inst_req_0); -- 
    convolve_cp_element_group_469: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_469"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(471);
      gj_convolve_cp_element_group_469 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(469), clk => clk, reset => reset); --
    end block;
    -- CP-element group 470:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 470: predecessors 
    -- CP-element group 470: 	26 
    -- CP-element group 470: marked-predecessors 
    -- CP-element group 470: 	472 
    -- CP-element group 470: 	524 
    -- CP-element group 470: successors 
    -- CP-element group 470: 	472 
    -- CP-element group 470:  members (3) 
      -- CP-element group 470: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Update/$entry
      -- CP-element group 470: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Update/cr
      -- CP-element group 470: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_update_start_
      -- 
    cr_6237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(470), ack => slice_2445_inst_req_1); -- 
    convolve_cp_element_group_470: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_470"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(472) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_470 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(470), clk => clk, reset => reset); --
    end block;
    -- CP-element group 471:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 471: predecessors 
    -- CP-element group 471: 	469 
    -- CP-element group 471: successors 
    -- CP-element group 471: marked-successors 
    -- CP-element group 471: 	354 
    -- CP-element group 471: 	469 
    -- CP-element group 471: 	366 
    -- CP-element group 471: 	378 
    -- CP-element group 471:  members (3) 
      -- CP-element group 471: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Sample/$exit
      -- CP-element group 471: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Sample/ra
      -- CP-element group 471: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_sample_completed_
      -- 
    ra_6233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 471_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2445_inst_ack_0, ack => convolve_CP_4675_elements(471)); -- 
    -- CP-element group 472:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 472: predecessors 
    -- CP-element group 472: 	470 
    -- CP-element group 472: successors 
    -- CP-element group 472: 	522 
    -- CP-element group 472: marked-successors 
    -- CP-element group 472: 	48 
    -- CP-element group 472: 	470 
    -- CP-element group 472: 	29 
    -- CP-element group 472:  members (3) 
      -- CP-element group 472: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Update/$exit
      -- CP-element group 472: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_Update/ca
      -- CP-element group 472: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2445_update_completed_
      -- 
    ca_6238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 472_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2445_inst_ack_1, ack => convolve_CP_4675_elements(472)); -- 
    -- CP-element group 473:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 473: predecessors 
    -- CP-element group 473: 	356 
    -- CP-element group 473: 	368 
    -- CP-element group 473: 	380 
    -- CP-element group 473: marked-predecessors 
    -- CP-element group 473: 	475 
    -- CP-element group 473: successors 
    -- CP-element group 473: 	475 
    -- CP-element group 473:  members (3) 
      -- CP-element group 473: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Sample/$entry
      -- CP-element group 473: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Sample/rr
      -- CP-element group 473: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_sample_start_
      -- 
    rr_6246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(473), ack => slice_2449_inst_req_0); -- 
    convolve_cp_element_group_473: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_473"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(475);
      gj_convolve_cp_element_group_473 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(473), clk => clk, reset => reset); --
    end block;
    -- CP-element group 474:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 474: predecessors 
    -- CP-element group 474: 	26 
    -- CP-element group 474: marked-predecessors 
    -- CP-element group 474: 	476 
    -- CP-element group 474: 	524 
    -- CP-element group 474: successors 
    -- CP-element group 474: 	476 
    -- CP-element group 474:  members (3) 
      -- CP-element group 474: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_update_start_
      -- CP-element group 474: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Update/cr
      -- CP-element group 474: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Update/$entry
      -- 
    cr_6251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(474), ack => slice_2449_inst_req_1); -- 
    convolve_cp_element_group_474: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_474"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(476) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_474 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(474), clk => clk, reset => reset); --
    end block;
    -- CP-element group 475:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 475: predecessors 
    -- CP-element group 475: 	473 
    -- CP-element group 475: successors 
    -- CP-element group 475: marked-successors 
    -- CP-element group 475: 	473 
    -- CP-element group 475: 	354 
    -- CP-element group 475: 	366 
    -- CP-element group 475: 	378 
    -- CP-element group 475:  members (3) 
      -- CP-element group 475: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Sample/ra
      -- CP-element group 475: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_sample_completed_
      -- CP-element group 475: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Sample/$exit
      -- 
    ra_6247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 475_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2449_inst_ack_0, ack => convolve_CP_4675_elements(475)); -- 
    -- CP-element group 476:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 476: predecessors 
    -- CP-element group 476: 	474 
    -- CP-element group 476: successors 
    -- CP-element group 476: 	522 
    -- CP-element group 476: marked-successors 
    -- CP-element group 476: 	474 
    -- CP-element group 476: 	48 
    -- CP-element group 476: 	29 
    -- CP-element group 476:  members (3) 
      -- CP-element group 476: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_update_completed_
      -- CP-element group 476: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Update/ca
      -- CP-element group 476: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/slice_2449_Update/$exit
      -- 
    ca_6252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 476_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_2449_inst_ack_1, ack => convolve_CP_4675_elements(476)); -- 
    -- CP-element group 477:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 477: predecessors 
    -- CP-element group 477: 	34 
    -- CP-element group 477: marked-predecessors 
    -- CP-element group 477: 	479 
    -- CP-element group 477: successors 
    -- CP-element group 477: 	479 
    -- CP-element group 477:  members (3) 
      -- CP-element group 477: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Sample/$entry
      -- CP-element group 477: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Sample/req
      -- CP-element group 477: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_sample_start_
      -- 
    req_6260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(477), ack => W_acc1_2884_delayed_2_0_2937_inst_req_0); -- 
    convolve_cp_element_group_477: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_477"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(34) & convolve_CP_4675_elements(479);
      gj_convolve_cp_element_group_477 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(477), clk => clk, reset => reset); --
    end block;
    -- CP-element group 478:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 478: predecessors 
    -- CP-element group 478: 	26 
    -- CP-element group 478: marked-predecessors 
    -- CP-element group 478: 	480 
    -- CP-element group 478: 	524 
    -- CP-element group 478: successors 
    -- CP-element group 478: 	480 
    -- CP-element group 478:  members (3) 
      -- CP-element group 478: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_update_start_
      -- CP-element group 478: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Update/$entry
      -- CP-element group 478: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Update/req
      -- 
    req_6265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(478), ack => W_acc1_2884_delayed_2_0_2937_inst_req_1); -- 
    convolve_cp_element_group_478: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_478"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(480) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_478 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(478), clk => clk, reset => reset); --
    end block;
    -- CP-element group 479:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 479: predecessors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: successors 
    -- CP-element group 479: marked-successors 
    -- CP-element group 479: 	477 
    -- CP-element group 479: 	30 
    -- CP-element group 479:  members (3) 
      -- CP-element group 479: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_sample_completed_
      -- CP-element group 479: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Sample/$exit
      -- CP-element group 479: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Sample/ack
      -- 
    ack_6261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 479_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2884_delayed_2_0_2937_inst_ack_0, ack => convolve_CP_4675_elements(479)); -- 
    -- CP-element group 480:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 480: predecessors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: successors 
    -- CP-element group 480: 	522 
    -- CP-element group 480: marked-successors 
    -- CP-element group 480: 	478 
    -- CP-element group 480: 	29 
    -- CP-element group 480:  members (3) 
      -- CP-element group 480: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_update_completed_
      -- CP-element group 480: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Update/ack
      -- CP-element group 480: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2939_Update/$exit
      -- 
    ack_6266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 480_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc1_2884_delayed_2_0_2937_inst_ack_1, ack => convolve_CP_4675_elements(480)); -- 
    -- CP-element group 481:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 481: predecessors 
    -- CP-element group 481: 	53 
    -- CP-element group 481: marked-predecessors 
    -- CP-element group 481: 	483 
    -- CP-element group 481: successors 
    -- CP-element group 481: 	483 
    -- CP-element group 481:  members (3) 
      -- CP-element group 481: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Sample/$entry
      -- CP-element group 481: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Sample/req
      -- CP-element group 481: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_sample_start_
      -- 
    req_6274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(481), ack => W_acc2_2893_delayed_2_0_2949_inst_req_0); -- 
    convolve_cp_element_group_481: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_481"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(53) & convolve_CP_4675_elements(483);
      gj_convolve_cp_element_group_481 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(481), clk => clk, reset => reset); --
    end block;
    -- CP-element group 482:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 482: predecessors 
    -- CP-element group 482: 	26 
    -- CP-element group 482: marked-predecessors 
    -- CP-element group 482: 	524 
    -- CP-element group 482: 	484 
    -- CP-element group 482: successors 
    -- CP-element group 482: 	484 
    -- CP-element group 482:  members (3) 
      -- CP-element group 482: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_update_start_
      -- CP-element group 482: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Update/$entry
      -- CP-element group 482: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Update/req
      -- 
    req_6279_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6279_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(482), ack => W_acc2_2893_delayed_2_0_2949_inst_req_1); -- 
    convolve_cp_element_group_482: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_482"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(484);
      gj_convolve_cp_element_group_482 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(482), clk => clk, reset => reset); --
    end block;
    -- CP-element group 483:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 483: predecessors 
    -- CP-element group 483: 	481 
    -- CP-element group 483: successors 
    -- CP-element group 483: marked-successors 
    -- CP-element group 483: 	481 
    -- CP-element group 483: 	49 
    -- CP-element group 483:  members (3) 
      -- CP-element group 483: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_sample_completed_
      -- CP-element group 483: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Sample/$exit
      -- CP-element group 483: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Sample/ack
      -- 
    ack_6275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 483_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2893_delayed_2_0_2949_inst_ack_0, ack => convolve_CP_4675_elements(483)); -- 
    -- CP-element group 484:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 484: predecessors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: successors 
    -- CP-element group 484: 	522 
    -- CP-element group 484: marked-successors 
    -- CP-element group 484: 	482 
    -- CP-element group 484: 	48 
    -- CP-element group 484:  members (3) 
      -- CP-element group 484: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_update_completed_
      -- CP-element group 484: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Update/$exit
      -- CP-element group 484: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_2951_Update/ack
      -- 
    ack_6280_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 484_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_acc2_2893_delayed_2_0_2949_inst_ack_1, ack => convolve_CP_4675_elements(484)); -- 
    -- CP-element group 485:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 485: predecessors 
    -- CP-element group 485: 	23 
    -- CP-element group 485: marked-predecessors 
    -- CP-element group 485: 	487 
    -- CP-element group 485: successors 
    -- CP-element group 485: 	487 
    -- CP-element group 485:  members (3) 
      -- CP-element group 485: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_sample_start_
      -- CP-element group 485: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Sample/rr
      -- CP-element group 485: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Sample/$entry
      -- 
    rr_6288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(485), ack => SUB_u16_u16_2986_inst_req_0); -- 
    convolve_cp_element_group_485: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_485"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(23) & convolve_CP_4675_elements(487);
      gj_convolve_cp_element_group_485 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(485), clk => clk, reset => reset); --
    end block;
    -- CP-element group 486:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 486: predecessors 
    -- CP-element group 486: marked-predecessors 
    -- CP-element group 486: 	498 
    -- CP-element group 486: 	505 
    -- CP-element group 486: 	491 
    -- CP-element group 486: 	488 
    -- CP-element group 486: successors 
    -- CP-element group 486: 	488 
    -- CP-element group 486:  members (3) 
      -- CP-element group 486: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Update/cr
      -- CP-element group 486: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Update/$entry
      -- CP-element group 486: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_update_start_
      -- 
    cr_6293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(486), ack => SUB_u16_u16_2986_inst_req_1); -- 
    convolve_cp_element_group_486: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_486"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(498) & convolve_CP_4675_elements(505) & convolve_CP_4675_elements(491) & convolve_CP_4675_elements(488);
      gj_convolve_cp_element_group_486 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(486), clk => clk, reset => reset); --
    end block;
    -- CP-element group 487:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 487: predecessors 
    -- CP-element group 487: 	485 
    -- CP-element group 487: successors 
    -- CP-element group 487: marked-successors 
    -- CP-element group 487: 	485 
    -- CP-element group 487:  members (3) 
      -- CP-element group 487: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_sample_completed_
      -- CP-element group 487: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Sample/ra
      -- CP-element group 487: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Sample/$exit
      -- 
    ra_6289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 487_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2986_inst_ack_0, ack => convolve_CP_4675_elements(487)); -- 
    -- CP-element group 488:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 488: predecessors 
    -- CP-element group 488: 	486 
    -- CP-element group 488: successors 
    -- CP-element group 488: 	24 
    -- CP-element group 488: 	496 
    -- CP-element group 488: 	503 
    -- CP-element group 488: 	489 
    -- CP-element group 488: marked-successors 
    -- CP-element group 488: 	486 
    -- CP-element group 488:  members (3) 
      -- CP-element group 488: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Update/$exit
      -- CP-element group 488: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_Update/ca
      -- CP-element group 488: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/SUB_u16_u16_2986_update_completed_
      -- 
    ca_6294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 488_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_2986_inst_ack_1, ack => convolve_CP_4675_elements(488)); -- 
    -- CP-element group 489:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 489: predecessors 
    -- CP-element group 489: 	72 
    -- CP-element group 489: 	91 
    -- CP-element group 489: 	488 
    -- CP-element group 489: marked-predecessors 
    -- CP-element group 489: 	491 
    -- CP-element group 489: successors 
    -- CP-element group 489: 	491 
    -- CP-element group 489:  members (3) 
      -- CP-element group 489: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_sample_start_
      -- CP-element group 489: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Sample/$entry
      -- CP-element group 489: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Sample/req
      -- 
    req_6302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(489), ack => W_store_kernel_2941_delayed_1_0_3004_inst_req_0); -- 
    convolve_cp_element_group_489: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_489"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(488) & convolve_CP_4675_elements(491);
      gj_convolve_cp_element_group_489 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(489), clk => clk, reset => reset); --
    end block;
    -- CP-element group 490:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 490: predecessors 
    -- CP-element group 490: marked-predecessors 
    -- CP-element group 490: 	492 
    -- CP-element group 490: 	494 
    -- CP-element group 490: successors 
    -- CP-element group 490: 	492 
    -- CP-element group 490:  members (3) 
      -- CP-element group 490: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Update/$entry
      -- CP-element group 490: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_update_start_
      -- CP-element group 490: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Update/req
      -- 
    req_6307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(490), ack => W_store_kernel_2941_delayed_1_0_3004_inst_req_1); -- 
    convolve_cp_element_group_490: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_490"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(492) & convolve_CP_4675_elements(494);
      gj_convolve_cp_element_group_490 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(490), clk => clk, reset => reset); --
    end block;
    -- CP-element group 491:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 491: predecessors 
    -- CP-element group 491: 	489 
    -- CP-element group 491: successors 
    -- CP-element group 491: marked-successors 
    -- CP-element group 491: 	87 
    -- CP-element group 491: 	68 
    -- CP-element group 491: 	486 
    -- CP-element group 491: 	489 
    -- CP-element group 491:  members (3) 
      -- CP-element group 491: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_sample_completed_
      -- CP-element group 491: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Sample/$exit
      -- CP-element group 491: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Sample/ack
      -- 
    ack_6303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 491_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2941_delayed_1_0_3004_inst_ack_0, ack => convolve_CP_4675_elements(491)); -- 
    -- CP-element group 492:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 492: predecessors 
    -- CP-element group 492: 	490 
    -- CP-element group 492: successors 
    -- CP-element group 492: 	493 
    -- CP-element group 492: marked-successors 
    -- CP-element group 492: 	490 
    -- CP-element group 492:  members (3) 
      -- CP-element group 492: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Update/$exit
      -- CP-element group 492: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_update_completed_
      -- CP-element group 492: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3006_Update/ack
      -- 
    ack_6308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 492_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2941_delayed_1_0_3004_inst_ack_1, ack => convolve_CP_4675_elements(492)); -- 
    -- CP-element group 493:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 493: predecessors 
    -- CP-element group 493: 	348 
    -- CP-element group 493: 	360 
    -- CP-element group 493: 	372 
    -- CP-element group 493: 	492 
    -- CP-element group 493: marked-predecessors 
    -- CP-element group 493: 	495 
    -- CP-element group 493: successors 
    -- CP-element group 493: 	494 
    -- CP-element group 493:  members (3) 
      -- CP-element group 493: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Sample/$entry
      -- CP-element group 493: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Sample/req
      -- CP-element group 493: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_sample_start_
      -- 
    req_6316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(493), ack => WPIPE_xxconvolvexxconv_k1_3008_inst_req_0); -- 
    convolve_cp_element_group_493: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_493"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(348) & convolve_CP_4675_elements(360) & convolve_CP_4675_elements(372) & convolve_CP_4675_elements(492) & convolve_CP_4675_elements(495);
      gj_convolve_cp_element_group_493 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(493), clk => clk, reset => reset); --
    end block;
    -- CP-element group 494:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 494: predecessors 
    -- CP-element group 494: 	493 
    -- CP-element group 494: successors 
    -- CP-element group 494: 	495 
    -- CP-element group 494: marked-successors 
    -- CP-element group 494: 	346 
    -- CP-element group 494: 	358 
    -- CP-element group 494: 	370 
    -- CP-element group 494: 	490 
    -- CP-element group 494:  members (6) 
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Sample/ack
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Sample/$exit
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_update_start_
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Update/$entry
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_sample_completed_
      -- CP-element group 494: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Update/req
      -- 
    ack_6317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 494_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_3008_inst_ack_0, ack => convolve_CP_4675_elements(494)); -- 
    req_6321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(494), ack => WPIPE_xxconvolvexxconv_k1_3008_inst_req_1); -- 
    -- CP-element group 495:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 495: predecessors 
    -- CP-element group 495: 	494 
    -- CP-element group 495: successors 
    -- CP-element group 495: 	530 
    -- CP-element group 495: marked-successors 
    -- CP-element group 495: 	493 
    -- CP-element group 495:  members (3) 
      -- CP-element group 495: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Update/ack
      -- CP-element group 495: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_update_completed_
      -- CP-element group 495: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k1_3008_Update/$exit
      -- 
    ack_6322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 495_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k1_3008_inst_ack_1, ack => convolve_CP_4675_elements(495)); -- 
    -- CP-element group 496:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 496: predecessors 
    -- CP-element group 496: 	72 
    -- CP-element group 496: 	91 
    -- CP-element group 496: 	488 
    -- CP-element group 496: marked-predecessors 
    -- CP-element group 496: 	498 
    -- CP-element group 496: successors 
    -- CP-element group 496: 	498 
    -- CP-element group 496:  members (3) 
      -- CP-element group 496: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_sample_start_
      -- CP-element group 496: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Sample/$entry
      -- CP-element group 496: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Sample/req
      -- 
    req_6330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(496), ack => W_store_kernel_2945_delayed_1_0_3011_inst_req_0); -- 
    convolve_cp_element_group_496: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_496"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(488) & convolve_CP_4675_elements(498);
      gj_convolve_cp_element_group_496 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(496), clk => clk, reset => reset); --
    end block;
    -- CP-element group 497:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 497: predecessors 
    -- CP-element group 497: marked-predecessors 
    -- CP-element group 497: 	499 
    -- CP-element group 497: 	501 
    -- CP-element group 497: successors 
    -- CP-element group 497: 	499 
    -- CP-element group 497:  members (3) 
      -- CP-element group 497: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_update_start_
      -- CP-element group 497: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Update/$entry
      -- CP-element group 497: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Update/req
      -- 
    req_6335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(497), ack => W_store_kernel_2945_delayed_1_0_3011_inst_req_1); -- 
    convolve_cp_element_group_497: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_497"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(499) & convolve_CP_4675_elements(501);
      gj_convolve_cp_element_group_497 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(497), clk => clk, reset => reset); --
    end block;
    -- CP-element group 498:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 498: predecessors 
    -- CP-element group 498: 	496 
    -- CP-element group 498: successors 
    -- CP-element group 498: marked-successors 
    -- CP-element group 498: 	496 
    -- CP-element group 498: 	87 
    -- CP-element group 498: 	68 
    -- CP-element group 498: 	486 
    -- CP-element group 498:  members (3) 
      -- CP-element group 498: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_sample_completed_
      -- CP-element group 498: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Sample/$exit
      -- CP-element group 498: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Sample/ack
      -- 
    ack_6331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 498_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2945_delayed_1_0_3011_inst_ack_0, ack => convolve_CP_4675_elements(498)); -- 
    -- CP-element group 499:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 499: predecessors 
    -- CP-element group 499: 	497 
    -- CP-element group 499: successors 
    -- CP-element group 499: 	500 
    -- CP-element group 499: marked-successors 
    -- CP-element group 499: 	497 
    -- CP-element group 499:  members (3) 
      -- CP-element group 499: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_update_completed_
      -- CP-element group 499: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Update/$exit
      -- CP-element group 499: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3013_Update/ack
      -- 
    ack_6336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 499_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2945_delayed_1_0_3011_inst_ack_1, ack => convolve_CP_4675_elements(499)); -- 
    -- CP-element group 500:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 500: predecessors 
    -- CP-element group 500: 	352 
    -- CP-element group 500: 	499 
    -- CP-element group 500: 	364 
    -- CP-element group 500: 	376 
    -- CP-element group 500: marked-predecessors 
    -- CP-element group 500: 	502 
    -- CP-element group 500: successors 
    -- CP-element group 500: 	501 
    -- CP-element group 500:  members (3) 
      -- CP-element group 500: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_sample_start_
      -- CP-element group 500: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Sample/$entry
      -- CP-element group 500: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Sample/req
      -- 
    req_6344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(500), ack => WPIPE_xxconvolvexxconv_k2_3015_inst_req_0); -- 
    convolve_cp_element_group_500: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_500"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(352) & convolve_CP_4675_elements(499) & convolve_CP_4675_elements(364) & convolve_CP_4675_elements(376) & convolve_CP_4675_elements(502);
      gj_convolve_cp_element_group_500 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(500), clk => clk, reset => reset); --
    end block;
    -- CP-element group 501:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 501: predecessors 
    -- CP-element group 501: 	500 
    -- CP-element group 501: successors 
    -- CP-element group 501: 	502 
    -- CP-element group 501: marked-successors 
    -- CP-element group 501: 	362 
    -- CP-element group 501: 	350 
    -- CP-element group 501: 	374 
    -- CP-element group 501: 	497 
    -- CP-element group 501:  members (6) 
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_sample_completed_
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_update_start_
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Sample/$exit
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Sample/ack
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Update/$entry
      -- CP-element group 501: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Update/req
      -- 
    ack_6345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 501_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_3015_inst_ack_0, ack => convolve_CP_4675_elements(501)); -- 
    req_6349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(501), ack => WPIPE_xxconvolvexxconv_k2_3015_inst_req_1); -- 
    -- CP-element group 502:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 502: predecessors 
    -- CP-element group 502: 	501 
    -- CP-element group 502: successors 
    -- CP-element group 502: 	530 
    -- CP-element group 502: marked-successors 
    -- CP-element group 502: 	500 
    -- CP-element group 502:  members (3) 
      -- CP-element group 502: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_update_completed_
      -- CP-element group 502: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Update/$exit
      -- CP-element group 502: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k2_3015_Update/ack
      -- 
    ack_6350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 502_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k2_3015_inst_ack_1, ack => convolve_CP_4675_elements(502)); -- 
    -- CP-element group 503:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 503: predecessors 
    -- CP-element group 503: 	72 
    -- CP-element group 503: 	91 
    -- CP-element group 503: 	488 
    -- CP-element group 503: marked-predecessors 
    -- CP-element group 503: 	505 
    -- CP-element group 503: successors 
    -- CP-element group 503: 	505 
    -- CP-element group 503:  members (3) 
      -- CP-element group 503: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_sample_start_
      -- CP-element group 503: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Sample/$entry
      -- CP-element group 503: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Sample/req
      -- 
    req_6358_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6358_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(503), ack => W_store_kernel_2949_delayed_1_0_3018_inst_req_0); -- 
    convolve_cp_element_group_503: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_503"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(72) & convolve_CP_4675_elements(91) & convolve_CP_4675_elements(488) & convolve_CP_4675_elements(505);
      gj_convolve_cp_element_group_503 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(503), clk => clk, reset => reset); --
    end block;
    -- CP-element group 504:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 504: predecessors 
    -- CP-element group 504: marked-predecessors 
    -- CP-element group 504: 	506 
    -- CP-element group 504: 	508 
    -- CP-element group 504: successors 
    -- CP-element group 504: 	506 
    -- CP-element group 504:  members (3) 
      -- CP-element group 504: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_update_start_
      -- CP-element group 504: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Update/$entry
      -- CP-element group 504: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Update/req
      -- 
    req_6363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(504), ack => W_store_kernel_2949_delayed_1_0_3018_inst_req_1); -- 
    convolve_cp_element_group_504: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_504"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(506) & convolve_CP_4675_elements(508);
      gj_convolve_cp_element_group_504 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(504), clk => clk, reset => reset); --
    end block;
    -- CP-element group 505:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 505: predecessors 
    -- CP-element group 505: 	503 
    -- CP-element group 505: successors 
    -- CP-element group 505: marked-successors 
    -- CP-element group 505: 	87 
    -- CP-element group 505: 	68 
    -- CP-element group 505: 	503 
    -- CP-element group 505: 	486 
    -- CP-element group 505:  members (3) 
      -- CP-element group 505: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_sample_completed_
      -- CP-element group 505: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Sample/$exit
      -- CP-element group 505: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Sample/ack
      -- 
    ack_6359_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 505_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2949_delayed_1_0_3018_inst_ack_0, ack => convolve_CP_4675_elements(505)); -- 
    -- CP-element group 506:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 506: predecessors 
    -- CP-element group 506: 	504 
    -- CP-element group 506: successors 
    -- CP-element group 506: 	507 
    -- CP-element group 506: marked-successors 
    -- CP-element group 506: 	504 
    -- CP-element group 506:  members (3) 
      -- CP-element group 506: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_update_completed_
      -- CP-element group 506: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Update/$exit
      -- CP-element group 506: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3020_Update/ack
      -- 
    ack_6364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 506_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_store_kernel_2949_delayed_1_0_3018_inst_ack_1, ack => convolve_CP_4675_elements(506)); -- 
    -- CP-element group 507:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 507: predecessors 
    -- CP-element group 507: 	356 
    -- CP-element group 507: 	368 
    -- CP-element group 507: 	506 
    -- CP-element group 507: 	380 
    -- CP-element group 507: marked-predecessors 
    -- CP-element group 507: 	509 
    -- CP-element group 507: successors 
    -- CP-element group 507: 	508 
    -- CP-element group 507:  members (3) 
      -- CP-element group 507: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_sample_start_
      -- CP-element group 507: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Sample/$entry
      -- CP-element group 507: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Sample/req
      -- 
    req_6372_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6372_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(507), ack => WPIPE_xxconvolvexxconv_k3_3022_inst_req_0); -- 
    convolve_cp_element_group_507: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_507"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(356) & convolve_CP_4675_elements(368) & convolve_CP_4675_elements(506) & convolve_CP_4675_elements(380) & convolve_CP_4675_elements(509);
      gj_convolve_cp_element_group_507 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(507), clk => clk, reset => reset); --
    end block;
    -- CP-element group 508:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 508: predecessors 
    -- CP-element group 508: 	507 
    -- CP-element group 508: successors 
    -- CP-element group 508: 	509 
    -- CP-element group 508: marked-successors 
    -- CP-element group 508: 	354 
    -- CP-element group 508: 	504 
    -- CP-element group 508: 	366 
    -- CP-element group 508: 	378 
    -- CP-element group 508:  members (6) 
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_sample_completed_
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_update_start_
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Sample/$exit
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Sample/ack
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Update/$entry
      -- CP-element group 508: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Update/req
      -- 
    ack_6373_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 508_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_3022_inst_ack_0, ack => convolve_CP_4675_elements(508)); -- 
    req_6377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(508), ack => WPIPE_xxconvolvexxconv_k3_3022_inst_req_1); -- 
    -- CP-element group 509:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 509: predecessors 
    -- CP-element group 509: 	508 
    -- CP-element group 509: successors 
    -- CP-element group 509: 	530 
    -- CP-element group 509: marked-successors 
    -- CP-element group 509: 	507 
    -- CP-element group 509:  members (3) 
      -- CP-element group 509: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_update_completed_
      -- CP-element group 509: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Update/$exit
      -- CP-element group 509: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_xxconvolvexxconv_k3_3022_Update/ack
      -- 
    ack_6378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 509_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_xxconvolvexxconv_k3_3022_inst_ack_1, ack => convolve_CP_4675_elements(509)); -- 
    -- CP-element group 510:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 510: predecessors 
    -- CP-element group 510: 	108 
    -- CP-element group 510: 	127 
    -- CP-element group 510: marked-predecessors 
    -- CP-element group 510: 	512 
    -- CP-element group 510: successors 
    -- CP-element group 510: 	512 
    -- CP-element group 510:  members (3) 
      -- CP-element group 510: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_sample_start_
      -- CP-element group 510: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Sample/$entry
      -- CP-element group 510: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Sample/req
      -- 
    req_6386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(510), ack => W_num_done_2992_delayed_2_0_3063_inst_req_0); -- 
    convolve_cp_element_group_510: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_510"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(127) & convolve_CP_4675_elements(512);
      gj_convolve_cp_element_group_510 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(510), clk => clk, reset => reset); --
    end block;
    -- CP-element group 511:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 511: predecessors 
    -- CP-element group 511: 	26 
    -- CP-element group 511: marked-predecessors 
    -- CP-element group 511: 	513 
    -- CP-element group 511: successors 
    -- CP-element group 511: 	513 
    -- CP-element group 511:  members (3) 
      -- CP-element group 511: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_update_start_
      -- CP-element group 511: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Update/$entry
      -- CP-element group 511: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Update/req
      -- 
    req_6391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(511), ack => W_num_done_2992_delayed_2_0_3063_inst_req_1); -- 
    convolve_cp_element_group_511: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_511"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(513);
      gj_convolve_cp_element_group_511 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(511), clk => clk, reset => reset); --
    end block;
    -- CP-element group 512:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 512: predecessors 
    -- CP-element group 512: 	510 
    -- CP-element group 512: successors 
    -- CP-element group 512: marked-successors 
    -- CP-element group 512: 	106 
    -- CP-element group 512: 	123 
    -- CP-element group 512: 	510 
    -- CP-element group 512:  members (3) 
      -- CP-element group 512: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_sample_completed_
      -- CP-element group 512: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Sample/$exit
      -- CP-element group 512: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Sample/ack
      -- 
    ack_6387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 512_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2992_delayed_2_0_3063_inst_ack_0, ack => convolve_CP_4675_elements(512)); -- 
    -- CP-element group 513:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 513: predecessors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: successors 
    -- CP-element group 513: 	530 
    -- CP-element group 513: marked-successors 
    -- CP-element group 513: 	511 
    -- CP-element group 513: 	29 
    -- CP-element group 513:  members (3) 
      -- CP-element group 513: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_update_completed_
      -- CP-element group 513: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Update/$exit
      -- CP-element group 513: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3065_Update/ack
      -- 
    ack_6392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 513_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2992_delayed_2_0_3063_inst_ack_1, ack => convolve_CP_4675_elements(513)); -- 
    -- CP-element group 514:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 514: predecessors 
    -- CP-element group 514: 	108 
    -- CP-element group 514: 	127 
    -- CP-element group 514: marked-predecessors 
    -- CP-element group 514: 	516 
    -- CP-element group 514: successors 
    -- CP-element group 514: 	516 
    -- CP-element group 514:  members (3) 
      -- CP-element group 514: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_sample_start_
      -- CP-element group 514: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Sample/$entry
      -- CP-element group 514: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Sample/req
      -- 
    req_6400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(514), ack => W_num_done_2998_delayed_2_0_3072_inst_req_0); -- 
    convolve_cp_element_group_514: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_514"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(127) & convolve_CP_4675_elements(516);
      gj_convolve_cp_element_group_514 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(514), clk => clk, reset => reset); --
    end block;
    -- CP-element group 515:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 515: predecessors 
    -- CP-element group 515: 	26 
    -- CP-element group 515: marked-predecessors 
    -- CP-element group 515: 	517 
    -- CP-element group 515: successors 
    -- CP-element group 515: 	517 
    -- CP-element group 515:  members (3) 
      -- CP-element group 515: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_update_start_
      -- CP-element group 515: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Update/$entry
      -- CP-element group 515: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Update/req
      -- 
    req_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(515), ack => W_num_done_2998_delayed_2_0_3072_inst_req_1); -- 
    convolve_cp_element_group_515: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_515"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(26) & convolve_CP_4675_elements(517);
      gj_convolve_cp_element_group_515 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(515), clk => clk, reset => reset); --
    end block;
    -- CP-element group 516:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 516: predecessors 
    -- CP-element group 516: 	514 
    -- CP-element group 516: successors 
    -- CP-element group 516: marked-successors 
    -- CP-element group 516: 	106 
    -- CP-element group 516: 	514 
    -- CP-element group 516: 	123 
    -- CP-element group 516:  members (3) 
      -- CP-element group 516: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_sample_completed_
      -- CP-element group 516: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Sample/$exit
      -- CP-element group 516: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Sample/ack
      -- 
    ack_6401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 516_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2998_delayed_2_0_3072_inst_ack_0, ack => convolve_CP_4675_elements(516)); -- 
    -- CP-element group 517:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 517: predecessors 
    -- CP-element group 517: 	515 
    -- CP-element group 517: successors 
    -- CP-element group 517: 	530 
    -- CP-element group 517: marked-successors 
    -- CP-element group 517: 	515 
    -- CP-element group 517: 	48 
    -- CP-element group 517:  members (3) 
      -- CP-element group 517: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_update_completed_
      -- CP-element group 517: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Update/$exit
      -- CP-element group 517: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3074_Update/ack
      -- 
    ack_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 517_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_2998_delayed_2_0_3072_inst_ack_1, ack => convolve_CP_4675_elements(517)); -- 
    -- CP-element group 518:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 518: predecessors 
    -- CP-element group 518: 	108 
    -- CP-element group 518: 	127 
    -- CP-element group 518: marked-predecessors 
    -- CP-element group 518: 	520 
    -- CP-element group 518: successors 
    -- CP-element group 518: 	520 
    -- CP-element group 518:  members (3) 
      -- CP-element group 518: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_sample_start_
      -- CP-element group 518: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Sample/$entry
      -- CP-element group 518: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Sample/req
      -- 
    req_6414_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6414_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(518), ack => W_num_done_3003_delayed_2_0_3081_inst_req_0); -- 
    convolve_cp_element_group_518: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_518"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(108) & convolve_CP_4675_elements(127) & convolve_CP_4675_elements(520);
      gj_convolve_cp_element_group_518 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(518), clk => clk, reset => reset); --
    end block;
    -- CP-element group 519:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 519: predecessors 
    -- CP-element group 519: marked-predecessors 
    -- CP-element group 519: 	521 
    -- CP-element group 519: 	524 
    -- CP-element group 519: 	527 
    -- CP-element group 519: successors 
    -- CP-element group 519: 	521 
    -- CP-element group 519:  members (3) 
      -- CP-element group 519: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_update_start_
      -- CP-element group 519: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Update/$entry
      -- CP-element group 519: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Update/req
      -- 
    req_6419_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6419_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(519), ack => W_num_done_3003_delayed_2_0_3081_inst_req_1); -- 
    convolve_cp_element_group_519: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_519"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(521) & convolve_CP_4675_elements(524) & convolve_CP_4675_elements(527);
      gj_convolve_cp_element_group_519 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(519), clk => clk, reset => reset); --
    end block;
    -- CP-element group 520:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 520: predecessors 
    -- CP-element group 520: 	518 
    -- CP-element group 520: successors 
    -- CP-element group 520: marked-successors 
    -- CP-element group 520: 	106 
    -- CP-element group 520: 	518 
    -- CP-element group 520: 	123 
    -- CP-element group 520:  members (3) 
      -- CP-element group 520: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_sample_completed_
      -- CP-element group 520: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Sample/$exit
      -- CP-element group 520: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Sample/ack
      -- 
    ack_6415_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 520_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3003_delayed_2_0_3081_inst_ack_0, ack => convolve_CP_4675_elements(520)); -- 
    -- CP-element group 521:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 521: predecessors 
    -- CP-element group 521: 	519 
    -- CP-element group 521: successors 
    -- CP-element group 521: 	522 
    -- CP-element group 521: 	526 
    -- CP-element group 521: marked-successors 
    -- CP-element group 521: 	519 
    -- CP-element group 521:  members (3) 
      -- CP-element group 521: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_update_completed_
      -- CP-element group 521: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Update/$exit
      -- CP-element group 521: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/assign_stmt_3083_Update/ack
      -- 
    ack_6420_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 521_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_num_done_3003_delayed_2_0_3081_inst_ack_1, ack => convolve_CP_4675_elements(521)); -- 
    -- CP-element group 522:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 522: predecessors 
    -- CP-element group 522: 	480 
    -- CP-element group 522: 	420 
    -- CP-element group 522: 	460 
    -- CP-element group 522: 	464 
    -- CP-element group 522: 	332 
    -- CP-element group 522: 	336 
    -- CP-element group 522: 	320 
    -- CP-element group 522: 	324 
    -- CP-element group 522: 	328 
    -- CP-element group 522: 	312 
    -- CP-element group 522: 	316 
    -- CP-element group 522: 	472 
    -- CP-element group 522: 	476 
    -- CP-element group 522: 	436 
    -- CP-element group 522: 	440 
    -- CP-element group 522: 	448 
    -- CP-element group 522: 	452 
    -- CP-element group 522: 	456 
    -- CP-element group 522: 	344 
    -- CP-element group 522: 	340 
    -- CP-element group 522: 	280 
    -- CP-element group 522: 	284 
    -- CP-element group 522: 	288 
    -- CP-element group 522: 	308 
    -- CP-element group 522: 	408 
    -- CP-element group 522: 	521 
    -- CP-element group 522: 	248 
    -- CP-element group 522: 	252 
    -- CP-element group 522: 	220 
    -- CP-element group 522: 	276 
    -- CP-element group 522: 	444 
    -- CP-element group 522: 	268 
    -- CP-element group 522: 	272 
    -- CP-element group 522: 	388 
    -- CP-element group 522: 	392 
    -- CP-element group 522: 	384 
    -- CP-element group 522: 	256 
    -- CP-element group 522: 	260 
    -- CP-element group 522: 	236 
    -- CP-element group 522: 	240 
    -- CP-element group 522: 	224 
    -- CP-element group 522: 	228 
    -- CP-element group 522: 	424 
    -- CP-element group 522: 	428 
    -- CP-element group 522: 	292 
    -- CP-element group 522: 	296 
    -- CP-element group 522: 	300 
    -- CP-element group 522: 	304 
    -- CP-element group 522: 	468 
    -- CP-element group 522: 	400 
    -- CP-element group 522: 	404 
    -- CP-element group 522: 	396 
    -- CP-element group 522: 	244 
    -- CP-element group 522: 	232 
    -- CP-element group 522: 	264 
    -- CP-element group 522: 	484 
    -- CP-element group 522: 	412 
    -- CP-element group 522: 	416 
    -- CP-element group 522: 	432 
    -- CP-element group 522: marked-predecessors 
    -- CP-element group 522: 	524 
    -- CP-element group 522: successors 
    -- CP-element group 522: 	524 
    -- CP-element group 522:  members (3) 
      -- CP-element group 522: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_sample_start_
      -- CP-element group 522: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Sample/$entry
      -- CP-element group 522: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Sample/rr
      -- 
    rr_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(522), ack => CONCAT_u8_u16_3090_inst_req_0); -- 
    convolve_cp_element_group_522: block -- 
      constant place_capacities: IntegerArray(0 to 59) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1,25 => 1,26 => 1,27 => 1,28 => 1,29 => 1,30 => 1,31 => 1,32 => 1,33 => 1,34 => 1,35 => 1,36 => 1,37 => 1,38 => 1,39 => 1,40 => 1,41 => 1,42 => 1,43 => 1,44 => 1,45 => 1,46 => 1,47 => 1,48 => 1,49 => 1,50 => 1,51 => 1,52 => 1,53 => 1,54 => 1,55 => 1,56 => 1,57 => 1,58 => 1,59 => 1);
      constant place_markings: IntegerArray(0 to 59)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0,41 => 0,42 => 0,43 => 0,44 => 0,45 => 0,46 => 0,47 => 0,48 => 0,49 => 0,50 => 0,51 => 0,52 => 0,53 => 0,54 => 0,55 => 0,56 => 0,57 => 0,58 => 0,59 => 1);
      constant place_delays: IntegerArray(0 to 59) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 0,25 => 0,26 => 0,27 => 0,28 => 0,29 => 0,30 => 0,31 => 0,32 => 0,33 => 0,34 => 0,35 => 0,36 => 0,37 => 0,38 => 0,39 => 0,40 => 0,41 => 0,42 => 0,43 => 0,44 => 0,45 => 0,46 => 0,47 => 0,48 => 0,49 => 0,50 => 0,51 => 0,52 => 0,53 => 0,54 => 0,55 => 0,56 => 0,57 => 0,58 => 0,59 => 1);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_522"; 
      signal preds: BooleanArray(1 to 60); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(480) & convolve_CP_4675_elements(420) & convolve_CP_4675_elements(460) & convolve_CP_4675_elements(464) & convolve_CP_4675_elements(332) & convolve_CP_4675_elements(336) & convolve_CP_4675_elements(320) & convolve_CP_4675_elements(324) & convolve_CP_4675_elements(328) & convolve_CP_4675_elements(312) & convolve_CP_4675_elements(316) & convolve_CP_4675_elements(472) & convolve_CP_4675_elements(476) & convolve_CP_4675_elements(436) & convolve_CP_4675_elements(440) & convolve_CP_4675_elements(448) & convolve_CP_4675_elements(452) & convolve_CP_4675_elements(456) & convolve_CP_4675_elements(344) & convolve_CP_4675_elements(340) & convolve_CP_4675_elements(280) & convolve_CP_4675_elements(284) & convolve_CP_4675_elements(288) & convolve_CP_4675_elements(308) & convolve_CP_4675_elements(408) & convolve_CP_4675_elements(521) & convolve_CP_4675_elements(248) & convolve_CP_4675_elements(252) & convolve_CP_4675_elements(220) & convolve_CP_4675_elements(276) & convolve_CP_4675_elements(444) & convolve_CP_4675_elements(268) & convolve_CP_4675_elements(272) & convolve_CP_4675_elements(388) & convolve_CP_4675_elements(392) & convolve_CP_4675_elements(384) & convolve_CP_4675_elements(256) & convolve_CP_4675_elements(260) & convolve_CP_4675_elements(236) & convolve_CP_4675_elements(240) & convolve_CP_4675_elements(224) & convolve_CP_4675_elements(228) & convolve_CP_4675_elements(424) & convolve_CP_4675_elements(428) & convolve_CP_4675_elements(292) & convolve_CP_4675_elements(296) & convolve_CP_4675_elements(300) & convolve_CP_4675_elements(304) & convolve_CP_4675_elements(468) & convolve_CP_4675_elements(400) & convolve_CP_4675_elements(404) & convolve_CP_4675_elements(396) & convolve_CP_4675_elements(244) & convolve_CP_4675_elements(232) & convolve_CP_4675_elements(264) & convolve_CP_4675_elements(484) & convolve_CP_4675_elements(412) & convolve_CP_4675_elements(416) & convolve_CP_4675_elements(432) & convolve_CP_4675_elements(524);
      gj_convolve_cp_element_group_522 : generic_join generic map(name => joinName, number_of_predecessors => 60, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(522), clk => clk, reset => reset); --
    end block;
    -- CP-element group 523:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 523: predecessors 
    -- CP-element group 523: marked-predecessors 
    -- CP-element group 523: 	525 
    -- CP-element group 523: 	527 
    -- CP-element group 523: successors 
    -- CP-element group 523: 	525 
    -- CP-element group 523:  members (3) 
      -- CP-element group 523: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_update_start_
      -- CP-element group 523: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Update/$entry
      -- CP-element group 523: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Update/cr
      -- 
    cr_6433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(523), ack => CONCAT_u8_u16_3090_inst_req_1); -- 
    convolve_cp_element_group_523: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_523"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(525) & convolve_CP_4675_elements(527);
      gj_convolve_cp_element_group_523 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(523), clk => clk, reset => reset); --
    end block;
    -- CP-element group 524:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 524: predecessors 
    -- CP-element group 524: 	522 
    -- CP-element group 524: successors 
    -- CP-element group 524: marked-successors 
    -- CP-element group 524: 	482 
    -- CP-element group 524: 	422 
    -- CP-element group 524: 	462 
    -- CP-element group 524: 	466 
    -- CP-element group 524: 	334 
    -- CP-element group 524: 	318 
    -- CP-element group 524: 	322 
    -- CP-element group 524: 	326 
    -- CP-element group 524: 	330 
    -- CP-element group 524: 	314 
    -- CP-element group 524: 	474 
    -- CP-element group 524: 	478 
    -- CP-element group 524: 	438 
    -- CP-element group 524: 	442 
    -- CP-element group 524: 	450 
    -- CP-element group 524: 	454 
    -- CP-element group 524: 	458 
    -- CP-element group 524: 	338 
    -- CP-element group 524: 	342 
    -- CP-element group 524: 	282 
    -- CP-element group 524: 	286 
    -- CP-element group 524: 	290 
    -- CP-element group 524: 	306 
    -- CP-element group 524: 	310 
    -- CP-element group 524: 	410 
    -- CP-element group 524: 	519 
    -- CP-element group 524: 	522 
    -- CP-element group 524: 	250 
    -- CP-element group 524: 	254 
    -- CP-element group 524: 	218 
    -- CP-element group 524: 	222 
    -- CP-element group 524: 	274 
    -- CP-element group 524: 	278 
    -- CP-element group 524: 	446 
    -- CP-element group 524: 	270 
    -- CP-element group 524: 	390 
    -- CP-element group 524: 	382 
    -- CP-element group 524: 	386 
    -- CP-element group 524: 	258 
    -- CP-element group 524: 	238 
    -- CP-element group 524: 	226 
    -- CP-element group 524: 	426 
    -- CP-element group 524: 	430 
    -- CP-element group 524: 	294 
    -- CP-element group 524: 	298 
    -- CP-element group 524: 	302 
    -- CP-element group 524: 	470 
    -- CP-element group 524: 	402 
    -- CP-element group 524: 	406 
    -- CP-element group 524: 	394 
    -- CP-element group 524: 	398 
    -- CP-element group 524: 	242 
    -- CP-element group 524: 	246 
    -- CP-element group 524: 	230 
    -- CP-element group 524: 	234 
    -- CP-element group 524: 	262 
    -- CP-element group 524: 	266 
    -- CP-element group 524: 	414 
    -- CP-element group 524: 	418 
    -- CP-element group 524: 	434 
    -- CP-element group 524:  members (3) 
      -- CP-element group 524: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_sample_completed_
      -- CP-element group 524: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Sample/$exit
      -- CP-element group 524: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Sample/ra
      -- 
    ra_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 524_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_3090_inst_ack_0, ack => convolve_CP_4675_elements(524)); -- 
    -- CP-element group 525:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 525: predecessors 
    -- CP-element group 525: 	523 
    -- CP-element group 525: successors 
    -- CP-element group 525: 	526 
    -- CP-element group 525: marked-successors 
    -- CP-element group 525: 	523 
    -- CP-element group 525:  members (3) 
      -- CP-element group 525: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_update_completed_
      -- CP-element group 525: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Update/$exit
      -- CP-element group 525: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/CONCAT_u8_u16_3090_Update/ca
      -- 
    ca_6434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 525_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u8_u16_3090_inst_ack_1, ack => convolve_CP_4675_elements(525)); -- 
    -- CP-element group 526:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 526: predecessors 
    -- CP-element group 526: 	521 
    -- CP-element group 526: 	525 
    -- CP-element group 526: marked-predecessors 
    -- CP-element group 526: 	528 
    -- CP-element group 526: successors 
    -- CP-element group 526: 	527 
    -- CP-element group 526:  members (3) 
      -- CP-element group 526: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_sample_start_
      -- CP-element group 526: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Sample/$entry
      -- CP-element group 526: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Sample/req
      -- 
    req_6442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(526), ack => WPIPE_output_pipe_3085_inst_req_0); -- 
    convolve_cp_element_group_526: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_526"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(521) & convolve_CP_4675_elements(525) & convolve_CP_4675_elements(528);
      gj_convolve_cp_element_group_526 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(526), clk => clk, reset => reset); --
    end block;
    -- CP-element group 527:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 527: predecessors 
    -- CP-element group 527: 	526 
    -- CP-element group 527: successors 
    -- CP-element group 527: 	528 
    -- CP-element group 527: marked-successors 
    -- CP-element group 527: 	519 
    -- CP-element group 527: 	523 
    -- CP-element group 527:  members (6) 
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_sample_completed_
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_update_start_
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Sample/$exit
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Sample/ack
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Update/$entry
      -- CP-element group 527: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Update/req
      -- 
    ack_6443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 527_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3085_inst_ack_0, ack => convolve_CP_4675_elements(527)); -- 
    req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(527), ack => WPIPE_output_pipe_3085_inst_req_1); -- 
    -- CP-element group 528:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 528: predecessors 
    -- CP-element group 528: 	527 
    -- CP-element group 528: successors 
    -- CP-element group 528: 	530 
    -- CP-element group 528: marked-successors 
    -- CP-element group 528: 	526 
    -- CP-element group 528:  members (3) 
      -- CP-element group 528: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_update_completed_
      -- CP-element group 528: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Update/$exit
      -- CP-element group 528: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/WPIPE_output_pipe_3085_Update/ack
      -- 
    ack_6448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 528_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_output_pipe_3085_inst_ack_1, ack => convolve_CP_4675_elements(528)); -- 
    -- CP-element group 529:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 529: predecessors 
    -- CP-element group 529: 	23 
    -- CP-element group 529: successors 
    -- CP-element group 529: 	24 
    -- CP-element group 529:  members (1) 
      -- CP-element group 529: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group convolve_CP_4675_elements(529) is a control-delay.
    cp_element_529_delay: control_delay_element  generic map(name => " 529_delay", delay_value => 1)  port map(req => convolve_CP_4675_elements(23), ack => convolve_CP_4675_elements(529), clk => clk, reset =>reset);
    -- CP-element group 530:  join  transition  bypass  pipeline-parent 
    -- CP-element group 530: predecessors 
    -- CP-element group 530: 	513 
    -- CP-element group 530: 	517 
    -- CP-element group 530: 	216 
    -- CP-element group 530: 	195 
    -- CP-element group 530: 	202 
    -- CP-element group 530: 	509 
    -- CP-element group 530: 	495 
    -- CP-element group 530: 	26 
    -- CP-element group 530: 	528 
    -- CP-element group 530: 	502 
    -- CP-element group 530: 	209 
    -- CP-element group 530: successors 
    -- CP-element group 530: 	20 
    -- CP-element group 530:  members (1) 
      -- CP-element group 530: 	 branch_block_stmt_1873/do_while_stmt_1890/do_while_stmt_1890_loop_body/$exit
      -- 
    convolve_cp_element_group_530: block -- 
      constant place_capacities: IntegerArray(0 to 10) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15,9 => 15,10 => 15);
      constant place_markings: IntegerArray(0 to 10)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant place_delays: IntegerArray(0 to 10) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0);
      constant joinName: string(1 to 29) := "convolve_cp_element_group_530"; 
      signal preds: BooleanArray(1 to 11); -- 
    begin -- 
      preds <= convolve_CP_4675_elements(513) & convolve_CP_4675_elements(517) & convolve_CP_4675_elements(216) & convolve_CP_4675_elements(195) & convolve_CP_4675_elements(202) & convolve_CP_4675_elements(509) & convolve_CP_4675_elements(495) & convolve_CP_4675_elements(26) & convolve_CP_4675_elements(528) & convolve_CP_4675_elements(502) & convolve_CP_4675_elements(209);
      gj_convolve_cp_element_group_530 : generic_join generic map(name => joinName, number_of_predecessors => 11, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convolve_CP_4675_elements(530), clk => clk, reset => reset); --
    end block;
    -- CP-element group 531:  transition  input  bypass  pipeline-parent 
    -- CP-element group 531: predecessors 
    -- CP-element group 531: 	19 
    -- CP-element group 531: successors 
    -- CP-element group 531:  members (2) 
      -- CP-element group 531: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_exit/$exit
      -- CP-element group 531: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_exit/ack
      -- 
    ack_6453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 531_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1890_branch_ack_0, ack => convolve_CP_4675_elements(531)); -- 
    -- CP-element group 532:  transition  input  bypass  pipeline-parent 
    -- CP-element group 532: predecessors 
    -- CP-element group 532: 	19 
    -- CP-element group 532: successors 
    -- CP-element group 532:  members (2) 
      -- CP-element group 532: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_taken/$exit
      -- CP-element group 532: 	 branch_block_stmt_1873/do_while_stmt_1890/loop_taken/ack
      -- 
    ack_6457_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 532_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1890_branch_ack_1, ack => convolve_CP_4675_elements(532)); -- 
    -- CP-element group 533:  transition  bypass  pipeline-parent 
    -- CP-element group 533: predecessors 
    -- CP-element group 533: 	17 
    -- CP-element group 533: successors 
    -- CP-element group 533: 	2 
    -- CP-element group 533:  members (1) 
      -- CP-element group 533: 	 branch_block_stmt_1873/do_while_stmt_1890/$exit
      -- 
    convolve_CP_4675_elements(533) <= convolve_CP_4675_elements(17);
    -- CP-element group 534:  transition  input  output  bypass 
    -- CP-element group 534: predecessors 
    -- CP-element group 534: 	2 
    -- CP-element group 534: successors 
    -- CP-element group 534: 	535 
    -- CP-element group 534:  members (6) 
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_sample_completed_
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_update_start_
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Sample/$exit
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Sample/ack
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Update/$entry
      -- CP-element group 534: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Update/req
      -- 
    ack_6470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 534_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3095_inst_ack_0, ack => convolve_CP_4675_elements(534)); -- 
    req_6474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(534), ack => WPIPE_input_done_pipe_3095_inst_req_1); -- 
    -- CP-element group 535:  transition  place  input  bypass 
    -- CP-element group 535: predecessors 
    -- CP-element group 535: 	534 
    -- CP-element group 535: successors 
    -- CP-element group 535: 	536 
    -- CP-element group 535:  members (8) 
      -- CP-element group 535: 	 branch_block_stmt_1873/assign_stmt_3097__exit__
      -- CP-element group 535: 	 branch_block_stmt_1873/loopback
      -- CP-element group 535: 	 branch_block_stmt_1873/assign_stmt_3097/$exit
      -- CP-element group 535: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_update_completed_
      -- CP-element group 535: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Update/$exit
      -- CP-element group 535: 	 branch_block_stmt_1873/assign_stmt_3097/WPIPE_input_done_pipe_3095_Update/ack
      -- CP-element group 535: 	 branch_block_stmt_1873/loopback_PhiReq/$entry
      -- CP-element group 535: 	 branch_block_stmt_1873/loopback_PhiReq/$exit
      -- 
    ack_6475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 535_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3095_inst_ack_1, ack => convolve_CP_4675_elements(535)); -- 
    -- CP-element group 536:  merge  fork  transition  place  output  bypass 
    -- CP-element group 536: predecessors 
    -- CP-element group 536: 	535 
    -- CP-element group 536: 	0 
    -- CP-element group 536: successors 
    -- CP-element group 536: 	3 
    -- CP-element group 536: 	6 
    -- CP-element group 536: 	14 
    -- CP-element group 536: 	11 
    -- CP-element group 536: 	10 
    -- CP-element group 536:  members (22) 
      -- CP-element group 536: 	 branch_block_stmt_1873/merge_stmt_1874__exit__
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889__entry__
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_num_out_pipe_1876_Sample/rr
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1878_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1883_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_update_start_
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_sample_start_
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Sample/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/RPIPE_size_pipe_1886_Sample/rr
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Update/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/assign_stmt_1879_to_assign_stmt_1889/SUB_u16_u16_1888_Update/cr
      -- CP-element group 536: 	 branch_block_stmt_1873/merge_stmt_1874_PhiReqMerge
      -- CP-element group 536: 	 branch_block_stmt_1873/merge_stmt_1874_PhiAck/$entry
      -- CP-element group 536: 	 branch_block_stmt_1873/merge_stmt_1874_PhiAck/$exit
      -- CP-element group 536: 	 branch_block_stmt_1873/merge_stmt_1874_PhiAck/dummy
      -- 
    rr_4706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(536), ack => RPIPE_num_out_pipe_1876_inst_req_0); -- 
    cr_4721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(536), ack => SUB_u16_u16_1878_inst_req_1); -- 
    cr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4749_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(536), ack => SUB_u16_u16_1883_inst_req_1); -- 
    rr_4762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(536), ack => RPIPE_size_pipe_1886_inst_req_0); -- 
    cr_4777_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4777_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convolve_CP_4675_elements(536), ack => SUB_u16_u16_1888_inst_req_1); -- 
    convolve_CP_4675_elements(536) <= OrReduce(convolve_CP_4675_elements(535) & convolve_CP_4675_elements(0));
    convolve_do_while_stmt_1890_terminator_6458: loop_terminator -- 
      generic map (name => " convolve_do_while_stmt_1890_terminator_6458", max_iterations_in_flight =>15) 
      port map(loop_body_exit => convolve_CP_4675_elements(20),loop_continue => convolve_CP_4675_elements(532),loop_terminate => convolve_CP_4675_elements(531),loop_back => convolve_CP_4675_elements(18),loop_exit => convolve_CP_4675_elements(17),clk => clk, reset => reset); -- 
    phi_stmt_1892_phi_seq_4842_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(37);
      convolve_CP_4675_elements(40)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(40);
      convolve_CP_4675_elements(41)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(42);
      convolve_CP_4675_elements(38) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(35);
      convolve_CP_4675_elements(44)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(46);
      convolve_CP_4675_elements(45)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(47);
      convolve_CP_4675_elements(36) <= phi_mux_reqs(1);
      phi_stmt_1892_phi_seq_4842 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1892_phi_seq_4842") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(31), 
          phi_sample_ack => convolve_CP_4675_elements(32), 
          phi_update_req => convolve_CP_4675_elements(33), 
          phi_update_ack => convolve_CP_4675_elements(34), 
          phi_mux_ack => convolve_CP_4675_elements(39), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1898_phi_seq_4886_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(56);
      convolve_CP_4675_elements(59)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(59);
      convolve_CP_4675_elements(60)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(61);
      convolve_CP_4675_elements(57) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(54);
      convolve_CP_4675_elements(63)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(65);
      convolve_CP_4675_elements(64)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(66);
      convolve_CP_4675_elements(55) <= phi_mux_reqs(1);
      phi_stmt_1898_phi_seq_4886 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1898_phi_seq_4886") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(50), 
          phi_sample_ack => convolve_CP_4675_elements(51), 
          phi_update_req => convolve_CP_4675_elements(52), 
          phi_update_ack => convolve_CP_4675_elements(53), 
          phi_mux_ack => convolve_CP_4675_elements(58), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1903_phi_seq_4930_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(75);
      convolve_CP_4675_elements(78)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(78);
      convolve_CP_4675_elements(79)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(80);
      convolve_CP_4675_elements(76) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(73);
      convolve_CP_4675_elements(82)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(84);
      convolve_CP_4675_elements(83)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(85);
      convolve_CP_4675_elements(74) <= phi_mux_reqs(1);
      phi_stmt_1903_phi_seq_4930 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1903_phi_seq_4930") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(69), 
          phi_sample_ack => convolve_CP_4675_elements(70), 
          phi_update_req => convolve_CP_4675_elements(71), 
          phi_update_ack => convolve_CP_4675_elements(72), 
          phi_mux_ack => convolve_CP_4675_elements(77), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1908_phi_seq_4974_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(94);
      convolve_CP_4675_elements(97)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(97);
      convolve_CP_4675_elements(98)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(99);
      convolve_CP_4675_elements(95) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(92);
      convolve_CP_4675_elements(101)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(103);
      convolve_CP_4675_elements(102)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(104);
      convolve_CP_4675_elements(93) <= phi_mux_reqs(1);
      phi_stmt_1908_phi_seq_4974 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1908_phi_seq_4974") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(88), 
          phi_sample_ack => convolve_CP_4675_elements(89), 
          phi_update_req => convolve_CP_4675_elements(90), 
          phi_update_ack => convolve_CP_4675_elements(91), 
          phi_mux_ack => convolve_CP_4675_elements(96), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1913_phi_seq_5018_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(111);
      convolve_CP_4675_elements(114)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(114);
      convolve_CP_4675_elements(115)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(116);
      convolve_CP_4675_elements(112) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(109);
      convolve_CP_4675_elements(118)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(120);
      convolve_CP_4675_elements(119)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(121);
      convolve_CP_4675_elements(110) <= phi_mux_reqs(1);
      phi_stmt_1913_phi_seq_5018 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1913_phi_seq_5018") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(25), 
          phi_sample_ack => convolve_CP_4675_elements(107), 
          phi_update_req => convolve_CP_4675_elements(27), 
          phi_update_ack => convolve_CP_4675_elements(108), 
          phi_mux_ack => convolve_CP_4675_elements(113), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1919_phi_seq_5062_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= convolve_CP_4675_elements(130);
      convolve_CP_4675_elements(133)<= src_sample_reqs(0);
      src_sample_acks(0)  <= convolve_CP_4675_elements(133);
      convolve_CP_4675_elements(134)<= src_update_reqs(0);
      src_update_acks(0)  <= convolve_CP_4675_elements(135);
      convolve_CP_4675_elements(131) <= phi_mux_reqs(0);
      triggers(1)  <= convolve_CP_4675_elements(128);
      convolve_CP_4675_elements(137)<= src_sample_reqs(1);
      src_sample_acks(1)  <= convolve_CP_4675_elements(139);
      convolve_CP_4675_elements(138)<= src_update_reqs(1);
      src_update_acks(1)  <= convolve_CP_4675_elements(140);
      convolve_CP_4675_elements(129) <= phi_mux_reqs(1);
      phi_stmt_1919_phi_seq_5062 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1919_phi_seq_5062") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => convolve_CP_4675_elements(124), 
          phi_sample_ack => convolve_CP_4675_elements(125), 
          phi_update_req => convolve_CP_4675_elements(126), 
          phi_update_ack => convolve_CP_4675_elements(127), 
          phi_mux_ack => convolve_CP_4675_elements(132), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_4794_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= convolve_CP_4675_elements(21);
        preds(1)  <= convolve_CP_4675_elements(22);
        entry_tmerge_4794 : transition_merge -- 
          generic map(name => " entry_tmerge_4794")
          port map (preds => preds, symbol_out => convolve_CP_4675_elements(23));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_i8_i8_2838_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2841_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2842_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2845_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2848_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2849_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2855_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2858_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2859_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2862_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2865_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2866_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2872_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2875_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2876_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2879_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2882_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2883_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2889_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2892_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2893_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2896_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2899_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2900_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2906_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2909_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2910_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2913_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2916_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2917_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2923_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2926_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2927_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2930_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2933_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2934_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2943_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2946_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2955_wire : std_logic_vector(7 downto 0);
    signal ADD_i8_i8_2958_wire : std_logic_vector(7 downto 0);
    signal ADD_u16_u16_3030_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3050_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3059_wire : std_logic_vector(15 downto 0);
    signal ADD_u2_u2_3039_wire : std_logic_vector(1 downto 0);
    signal AND_u1_u1_2996_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u8_u16_3090_wire : std_logic_vector(15 downto 0);
    signal EQ_u16_u1_1928_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2298_wire : std_logic_vector(0 downto 0);
    signal EQ_u16_u1_2301_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1931_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_2969_wire : std_logic_vector(0 downto 0);
    signal MUL_i8_i8_2550_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2556_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2562_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2568_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2574_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2580_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2586_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2592_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2598_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2604_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2610_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2616_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2622_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2628_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2634_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2640_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2646_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2652_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2658_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2664_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2670_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2676_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2682_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2688_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2694_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2700_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2706_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2712_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2718_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2724_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2730_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2736_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2742_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2748_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2754_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2760_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2766_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2772_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2778_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2784_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2790_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2796_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2802_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2808_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2814_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2820_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2826_wire : std_logic_vector(7 downto 0);
    signal MUL_i8_i8_2832_wire : std_logic_vector(7 downto 0);
    signal MUX_3040_wire : std_logic_vector(1 downto 0);
    signal MUX_3051_wire : std_logic_vector(15 downto 0);
    signal NOT_u1_u1_3094_wire : std_logic_vector(0 downto 0);
    signal RPIPE_num_out_pipe_1876_wire : std_logic_vector(15 downto 0);
    signal RPIPE_num_out_pipe_1881_wire : std_logic_vector(15 downto 0);
    signal RPIPE_size_pipe_1886_wire : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_2927_2927_delayed_1_0_2987 : std_logic_vector(15 downto 0);
    signal UGT_u2_u1_2008_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_2005_wire : std_logic_vector(0 downto 0);
    signal acc1_1892 : std_logic_vector(7 downto 0);
    signal acc1_2884_delayed_2_0_2939 : std_logic_vector(7 downto 0);
    signal acc2_1898 : std_logic_vector(7 downto 0);
    signal acc2_2893_delayed_2_0_2951 : std_logic_vector(7 downto 0);
    signal acc_val1_2948 : std_logic_vector(7 downto 0);
    signal acc_val2_2960 : std_logic_vector(7 downto 0);
    signal all_done_flag_3003 : std_logic_vector(0 downto 0);
    signal chl_1919 : std_logic_vector(15 downto 0);
    signal chl_done_2965 : std_logic_vector(0 downto 0);
    signal col_1908 : std_logic_vector(15 downto 0);
    signal col_done_2977 : std_logic_vector(0 downto 0);
    signal ir1_1_2042 : std_logic_vector(7 downto 0);
    signal ir1_2_2074 : std_logic_vector(7 downto 0);
    signal ir1_3_2106 : std_logic_vector(7 downto 0);
    signal ir1_4_2138 : std_logic_vector(7 downto 0);
    signal ir2_1_2046 : std_logic_vector(7 downto 0);
    signal ir2_2_2078 : std_logic_vector(7 downto 0);
    signal ir2_3_2110 : std_logic_vector(7 downto 0);
    signal ir2_4_2142 : std_logic_vector(7 downto 0);
    signal ir3_1_2050 : std_logic_vector(7 downto 0);
    signal ir3_2_2082 : std_logic_vector(7 downto 0);
    signal ir3_3_2114 : std_logic_vector(7 downto 0);
    signal ir3_4_2146 : std_logic_vector(7 downto 0);
    signal ir4_1_2054 : std_logic_vector(7 downto 0);
    signal ir4_2_2086 : std_logic_vector(7 downto 0);
    signal ir4_3_2118 : std_logic_vector(7 downto 0);
    signal ir4_4_2150 : std_logic_vector(7 downto 0);
    signal ir5_1_2058 : std_logic_vector(7 downto 0);
    signal ir5_2_2090 : std_logic_vector(7 downto 0);
    signal ir5_3_2122 : std_logic_vector(7 downto 0);
    signal ir5_4_2154 : std_logic_vector(7 downto 0);
    signal ir6_1_2062 : std_logic_vector(7 downto 0);
    signal ir6_2_2094 : std_logic_vector(7 downto 0);
    signal ir6_3_2126 : std_logic_vector(7 downto 0);
    signal ir6_4_2158 : std_logic_vector(7 downto 0);
    signal ir7_1_2066 : std_logic_vector(7 downto 0);
    signal ir7_2_2098 : std_logic_vector(7 downto 0);
    signal ir7_3_2130 : std_logic_vector(7 downto 0);
    signal ir7_4_2162 : std_logic_vector(7 downto 0);
    signal ir8_1_2070 : std_logic_vector(7 downto 0);
    signal ir8_2_2102 : std_logic_vector(7 downto 0);
    signal ir8_3_2134 : std_logic_vector(7 downto 0);
    signal ir8_4_2166 : std_logic_vector(7 downto 0);
    signal iread1_1974 : std_logic_vector(63 downto 0);
    signal iread2_1983 : std_logic_vector(63 downto 0);
    signal iread3_1992 : std_logic_vector(63 downto 0);
    signal iread4_2001 : std_logic_vector(63 downto 0);
    signal ival1_1_2170 : std_logic_vector(7 downto 0);
    signal ival1_2_2202 : std_logic_vector(7 downto 0);
    signal ival1_3_2234 : std_logic_vector(7 downto 0);
    signal ival1_4_2266 : std_logic_vector(7 downto 0);
    signal ival2_1_2174 : std_logic_vector(7 downto 0);
    signal ival2_2_2206 : std_logic_vector(7 downto 0);
    signal ival2_3_2238 : std_logic_vector(7 downto 0);
    signal ival2_4_2270 : std_logic_vector(7 downto 0);
    signal ival3_1_2178 : std_logic_vector(7 downto 0);
    signal ival3_2_2210 : std_logic_vector(7 downto 0);
    signal ival3_3_2242 : std_logic_vector(7 downto 0);
    signal ival3_4_2274 : std_logic_vector(7 downto 0);
    signal ival4_1_2182 : std_logic_vector(7 downto 0);
    signal ival4_2_2214 : std_logic_vector(7 downto 0);
    signal ival4_3_2246 : std_logic_vector(7 downto 0);
    signal ival4_4_2278 : std_logic_vector(7 downto 0);
    signal ival5_1_2186 : std_logic_vector(7 downto 0);
    signal ival5_2_2218 : std_logic_vector(7 downto 0);
    signal ival5_3_2250 : std_logic_vector(7 downto 0);
    signal ival5_4_2282 : std_logic_vector(7 downto 0);
    signal ival6_1_2190 : std_logic_vector(7 downto 0);
    signal ival6_2_2222 : std_logic_vector(7 downto 0);
    signal ival6_3_2254 : std_logic_vector(7 downto 0);
    signal ival6_4_2286 : std_logic_vector(7 downto 0);
    signal ival7_1_2194 : std_logic_vector(7 downto 0);
    signal ival7_2_2226 : std_logic_vector(7 downto 0);
    signal ival7_3_2258 : std_logic_vector(7 downto 0);
    signal ival7_4_2290 : std_logic_vector(7 downto 0);
    signal ival8_1_2198 : std_logic_vector(7 downto 0);
    signal ival8_2_2230 : std_logic_vector(7 downto 0);
    signal ival8_3_2262 : std_logic_vector(7 downto 0);
    signal ival8_4_2294 : std_logic_vector(7 downto 0);
    signal konst_1877_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1882_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1887_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1927_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1930_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2007_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2297_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2300_wire_constant : std_logic_vector(15 downto 0);
    signal konst_2968_wire_constant : std_logic_vector(1 downto 0);
    signal konst_2985_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3027_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3029_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3036_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3038_wire_constant : std_logic_vector(1 downto 0);
    signal konst_3047_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3049_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3058_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3068_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3077_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3096_wire_constant : std_logic_vector(7 downto 0);
    signal kr1_1_2358 : std_logic_vector(7 downto 0);
    signal kr1_2_2390 : std_logic_vector(7 downto 0);
    signal kr1_3_2422 : std_logic_vector(7 downto 0);
    signal kr2_1_2362 : std_logic_vector(7 downto 0);
    signal kr2_2_2394 : std_logic_vector(7 downto 0);
    signal kr2_3_2426 : std_logic_vector(7 downto 0);
    signal kr3_1_2366 : std_logic_vector(7 downto 0);
    signal kr3_2_2398 : std_logic_vector(7 downto 0);
    signal kr3_3_2430 : std_logic_vector(7 downto 0);
    signal kr4_1_2370 : std_logic_vector(7 downto 0);
    signal kr4_2_2402 : std_logic_vector(7 downto 0);
    signal kr4_3_2434 : std_logic_vector(7 downto 0);
    signal kr5_1_2374 : std_logic_vector(7 downto 0);
    signal kr5_2_2406 : std_logic_vector(7 downto 0);
    signal kr5_3_2438 : std_logic_vector(7 downto 0);
    signal kr6_1_2378 : std_logic_vector(7 downto 0);
    signal kr6_2_2410 : std_logic_vector(7 downto 0);
    signal kr6_3_2442 : std_logic_vector(7 downto 0);
    signal kr7_1_2382 : std_logic_vector(7 downto 0);
    signal kr7_2_2414 : std_logic_vector(7 downto 0);
    signal kr7_3_2446 : std_logic_vector(7 downto 0);
    signal kr8_1_2386 : std_logic_vector(7 downto 0);
    signal kr8_2_2418 : std_logic_vector(7 downto 0);
    signal kr8_3_2450 : std_logic_vector(7 downto 0);
    signal kread1_2336 : std_logic_vector(63 downto 0);
    signal kread2_2345 : std_logic_vector(63 downto 0);
    signal kread3_2354 : std_logic_vector(63 downto 0);
    signal kval1_1_2454 : std_logic_vector(7 downto 0);
    signal kval1_2_2486 : std_logic_vector(7 downto 0);
    signal kval1_3_2518 : std_logic_vector(7 downto 0);
    signal kval2_1_2458 : std_logic_vector(7 downto 0);
    signal kval2_2_2490 : std_logic_vector(7 downto 0);
    signal kval2_3_2522 : std_logic_vector(7 downto 0);
    signal kval3_1_2462 : std_logic_vector(7 downto 0);
    signal kval3_2_2494 : std_logic_vector(7 downto 0);
    signal kval3_3_2526 : std_logic_vector(7 downto 0);
    signal kval4_1_2466 : std_logic_vector(7 downto 0);
    signal kval4_2_2498 : std_logic_vector(7 downto 0);
    signal kval4_3_2530 : std_logic_vector(7 downto 0);
    signal kval5_1_2470 : std_logic_vector(7 downto 0);
    signal kval5_2_2502 : std_logic_vector(7 downto 0);
    signal kval5_3_2534 : std_logic_vector(7 downto 0);
    signal kval6_1_2474 : std_logic_vector(7 downto 0);
    signal kval6_2_2506 : std_logic_vector(7 downto 0);
    signal kval6_3_2538 : std_logic_vector(7 downto 0);
    signal kval7_1_2478 : std_logic_vector(7 downto 0);
    signal kval7_2_2510 : std_logic_vector(7 downto 0);
    signal kval7_3_2542 : std_logic_vector(7 downto 0);
    signal kval8_1_2482 : std_logic_vector(7 downto 0);
    signal kval8_2_2514 : std_logic_vector(7 downto 0);
    signal kval8_3_2546 : std_logic_vector(7 downto 0);
    signal mul_val1_1_2552 : std_logic_vector(7 downto 0);
    signal mul_val1_2_2600 : std_logic_vector(7 downto 0);
    signal mul_val1_3_2648 : std_logic_vector(7 downto 0);
    signal mul_val1_4_2696 : std_logic_vector(7 downto 0);
    signal mul_val1_5_2744 : std_logic_vector(7 downto 0);
    signal mul_val1_6_2792 : std_logic_vector(7 downto 0);
    signal mul_val2_1_2558 : std_logic_vector(7 downto 0);
    signal mul_val2_2_2606 : std_logic_vector(7 downto 0);
    signal mul_val2_3_2654 : std_logic_vector(7 downto 0);
    signal mul_val2_4_2702 : std_logic_vector(7 downto 0);
    signal mul_val2_5_2750 : std_logic_vector(7 downto 0);
    signal mul_val2_6_2798 : std_logic_vector(7 downto 0);
    signal mul_val3_1_2564 : std_logic_vector(7 downto 0);
    signal mul_val3_2_2612 : std_logic_vector(7 downto 0);
    signal mul_val3_3_2660 : std_logic_vector(7 downto 0);
    signal mul_val3_4_2708 : std_logic_vector(7 downto 0);
    signal mul_val3_5_2756 : std_logic_vector(7 downto 0);
    signal mul_val3_6_2804 : std_logic_vector(7 downto 0);
    signal mul_val4_1_2570 : std_logic_vector(7 downto 0);
    signal mul_val4_2_2618 : std_logic_vector(7 downto 0);
    signal mul_val4_3_2666 : std_logic_vector(7 downto 0);
    signal mul_val4_4_2714 : std_logic_vector(7 downto 0);
    signal mul_val4_5_2762 : std_logic_vector(7 downto 0);
    signal mul_val4_6_2810 : std_logic_vector(7 downto 0);
    signal mul_val5_1_2576 : std_logic_vector(7 downto 0);
    signal mul_val5_2_2624 : std_logic_vector(7 downto 0);
    signal mul_val5_3_2672 : std_logic_vector(7 downto 0);
    signal mul_val5_4_2720 : std_logic_vector(7 downto 0);
    signal mul_val5_5_2768 : std_logic_vector(7 downto 0);
    signal mul_val5_6_2816 : std_logic_vector(7 downto 0);
    signal mul_val6_1_2582 : std_logic_vector(7 downto 0);
    signal mul_val6_2_2630 : std_logic_vector(7 downto 0);
    signal mul_val6_3_2678 : std_logic_vector(7 downto 0);
    signal mul_val6_4_2726 : std_logic_vector(7 downto 0);
    signal mul_val6_5_2774 : std_logic_vector(7 downto 0);
    signal mul_val6_6_2822 : std_logic_vector(7 downto 0);
    signal mul_val7_1_2588 : std_logic_vector(7 downto 0);
    signal mul_val7_2_2636 : std_logic_vector(7 downto 0);
    signal mul_val7_3_2684 : std_logic_vector(7 downto 0);
    signal mul_val7_4_2732 : std_logic_vector(7 downto 0);
    signal mul_val7_5_2780 : std_logic_vector(7 downto 0);
    signal mul_val7_6_2828 : std_logic_vector(7 downto 0);
    signal mul_val8_1_2594 : std_logic_vector(7 downto 0);
    signal mul_val8_2_2642 : std_logic_vector(7 downto 0);
    signal mul_val8_3_2690 : std_logic_vector(7 downto 0);
    signal mul_val8_4_2738 : std_logic_vector(7 downto 0);
    signal mul_val8_5_2786 : std_logic_vector(7 downto 0);
    signal mul_val8_6_2834 : std_logic_vector(7 downto 0);
    signal n_chl_3032 : std_logic_vector(15 downto 0);
    signal n_chl_3032_1923_buffered : std_logic_vector(15 downto 0);
    signal n_col_3054 : std_logic_vector(15 downto 0);
    signal n_col_3054_1912_buffered : std_logic_vector(15 downto 0);
    signal n_num_3043 : std_logic_vector(1 downto 0);
    signal n_num_3043_1918_buffered : std_logic_vector(1 downto 0);
    signal n_row_3062 : std_logic_vector(15 downto 0);
    signal n_row_3062_1907_buffered : std_logic_vector(15 downto 0);
    signal nacc1_3071 : std_logic_vector(7 downto 0);
    signal nacc1_3071_1897_buffered : std_logic_vector(7 downto 0);
    signal nacc2_3080 : std_logic_vector(7 downto 0);
    signal nacc2_3080_1902_buffered : std_logic_vector(7 downto 0);
    signal num_1913 : std_logic_vector(1 downto 0);
    signal num_chl_1889 : std_logic_vector(15 downto 0);
    signal num_col_1884 : std_logic_vector(15 downto 0);
    signal num_done_2972 : std_logic_vector(0 downto 0);
    signal num_done_2992_delayed_2_0_3065 : std_logic_vector(0 downto 0);
    signal num_done_2998_delayed_2_0_3074 : std_logic_vector(0 downto 0);
    signal num_done_3003_delayed_2_0_3083 : std_logic_vector(0 downto 0);
    signal num_row_1879 : std_logic_vector(15 downto 0);
    signal out_done_flag_2992 : std_logic_vector(0 downto 0);
    signal read_ip_1933 : std_logic_vector(0 downto 0);
    signal read_ip_1946_delayed_1_0_1968 : std_logic_vector(0 downto 0);
    signal read_ip_1952_delayed_1_0_1977 : std_logic_vector(0 downto 0);
    signal read_ip_1958_delayed_1_0_1986 : std_logic_vector(0 downto 0);
    signal read_ip_1964_delayed_1_0_1995 : std_logic_vector(0 downto 0);
    signal read_k_2284_delayed_1_0_2330 : std_logic_vector(0 downto 0);
    signal read_k_2290_delayed_1_0_2339 : std_logic_vector(0 downto 0);
    signal read_k_2296_delayed_1_0_2348 : std_logic_vector(0 downto 0);
    signal read_k_2303 : std_logic_vector(0 downto 0);
    signal row_1903 : std_logic_vector(15 downto 0);
    signal row_done_2982 : std_logic_vector(0 downto 0);
    signal store_kernel_2941_delayed_1_0_3006 : std_logic_vector(0 downto 0);
    signal store_kernel_2945_delayed_1_0_3013 : std_logic_vector(0 downto 0);
    signal store_kernel_2949_delayed_1_0_3020 : std_logic_vector(0 downto 0);
    signal store_kernel_2998 : std_logic_vector(0 downto 0);
    signal t_acc_val1_2851 : std_logic_vector(7 downto 0);
    signal t_acc_val2_2868 : std_logic_vector(7 downto 0);
    signal t_acc_val3_2885 : std_logic_vector(7 downto 0);
    signal t_acc_val4_2902 : std_logic_vector(7 downto 0);
    signal t_acc_val5_2919 : std_logic_vector(7 downto 0);
    signal t_acc_val6_2936 : std_logic_vector(7 downto 0);
    signal temp1_1_1953 : std_logic_vector(63 downto 0);
    signal temp1_2_1957 : std_logic_vector(63 downto 0);
    signal temp1_3_1961 : std_logic_vector(63 downto 0);
    signal temp1_4_1965 : std_logic_vector(63 downto 0);
    signal temp2_1_1937 : std_logic_vector(63 downto 0);
    signal temp2_2_1941 : std_logic_vector(63 downto 0);
    signal temp2_3_1945 : std_logic_vector(63 downto 0);
    signal temp2_4_1949 : std_logic_vector(63 downto 0);
    signal tempk1_1_2307 : std_logic_vector(63 downto 0);
    signal tempk1_2_2311 : std_logic_vector(63 downto 0);
    signal tempk1_3_2315 : std_logic_vector(63 downto 0);
    signal tempk2_1_2319 : std_logic_vector(63 downto 0);
    signal tempk2_2_2323 : std_logic_vector(63 downto 0);
    signal tempk2_3_2327 : std_logic_vector(63 downto 0);
    signal type_cast_1896_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1901_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1906_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1911_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1917_wire_constant : std_logic_vector(1 downto 0);
    signal type_cast_1922_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3087_wire : std_logic_vector(7 downto 0);
    signal type_cast_3089_wire : std_logic_vector(7 downto 0);
    signal write_input_1978_delayed_1_0_2013 : std_logic_vector(0 downto 0);
    signal write_input_1982_delayed_1_0_2020 : std_logic_vector(0 downto 0);
    signal write_input_1986_delayed_1_0_2027 : std_logic_vector(0 downto 0);
    signal write_input_1990_delayed_1_0_2034 : std_logic_vector(0 downto 0);
    signal write_input_2010 : std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip1
    signal xxconvolvexxconv_ip1_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip2
    signal xxconvolvexxconv_ip2_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip3
    signal xxconvolvexxconv_ip3_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_ip4
    signal xxconvolvexxconv_ip4_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_ip4_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k1
    signal xxconvolvexxconv_k1_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k1_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k2
    signal xxconvolvexxconv_k2_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k2_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxconvolvexxconv_k3
    signal xxconvolvexxconv_k3_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxconvolvexxconv_k3_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1877_wire_constant <= "0000000000000001";
    konst_1882_wire_constant <= "0000000000000001";
    konst_1887_wire_constant <= "0000000000000001";
    konst_1927_wire_constant <= "0000000000000000";
    konst_1930_wire_constant <= "10";
    konst_2007_wire_constant <= "00";
    konst_2297_wire_constant <= "0000000000000000";
    konst_2300_wire_constant <= "0000000000000000";
    konst_2968_wire_constant <= "10";
    konst_2985_wire_constant <= "0000000000000001";
    konst_3027_wire_constant <= "0000000000000000";
    konst_3029_wire_constant <= "0000000000000001";
    konst_3036_wire_constant <= "00";
    konst_3038_wire_constant <= "01";
    konst_3047_wire_constant <= "0000000000000000";
    konst_3049_wire_constant <= "0000000000000001";
    konst_3058_wire_constant <= "0000000000000010";
    konst_3068_wire_constant <= "00000000";
    konst_3077_wire_constant <= "00000000";
    konst_3096_wire_constant <= "00000001";
    type_cast_1896_wire_constant <= "00000000";
    type_cast_1901_wire_constant <= "00000000";
    type_cast_1906_wire_constant <= "0000000000000000";
    type_cast_1911_wire_constant <= "0000000000000000";
    type_cast_1917_wire_constant <= "00";
    type_cast_1922_wire_constant <= "0000000000000000";
    phi_stmt_1892: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1896_wire_constant & nacc1_3071_1897_buffered;
      req <= phi_stmt_1892_req_0 & phi_stmt_1892_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1892",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1892_ack_0,
          idata => idata,
          odata => acc1_1892,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1892
    phi_stmt_1898: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1901_wire_constant & nacc2_3080_1902_buffered;
      req <= phi_stmt_1898_req_0 & phi_stmt_1898_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1898",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1898_ack_0,
          idata => idata,
          odata => acc2_1898,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1898
    phi_stmt_1903: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1906_wire_constant & n_row_3062_1907_buffered;
      req <= phi_stmt_1903_req_0 & phi_stmt_1903_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1903",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1903_ack_0,
          idata => idata,
          odata => row_1903,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1903
    phi_stmt_1908: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1911_wire_constant & n_col_3054_1912_buffered;
      req <= phi_stmt_1908_req_0 & phi_stmt_1908_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1908",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1908_ack_0,
          idata => idata,
          odata => col_1908,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1908
    phi_stmt_1913: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1917_wire_constant & n_num_3043_1918_buffered;
      req <= phi_stmt_1913_req_0 & phi_stmt_1913_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1913",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1913_ack_0,
          idata => idata,
          odata => num_1913,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1913
    phi_stmt_1919: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1922_wire_constant & n_chl_3032_1923_buffered;
      req <= phi_stmt_1919_req_0 & phi_stmt_1919_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1919",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1919_ack_0,
          idata => idata,
          odata => chl_1919,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1919
    -- flow-through select operator MUX_1973_inst
    iread1_1974 <= temp2_1_1937 when (read_ip_1946_delayed_1_0_1968(0) /=  '0') else temp1_1_1953;
    -- flow-through select operator MUX_1982_inst
    iread2_1983 <= temp2_2_1941 when (read_ip_1952_delayed_1_0_1977(0) /=  '0') else temp1_2_1957;
    -- flow-through select operator MUX_1991_inst
    iread3_1992 <= temp2_3_1945 when (read_ip_1958_delayed_1_0_1986(0) /=  '0') else temp1_3_1961;
    -- flow-through select operator MUX_2000_inst
    iread4_2001 <= temp2_4_1949 when (read_ip_1964_delayed_1_0_1995(0) /=  '0') else temp1_4_1965;
    -- flow-through select operator MUX_2335_inst
    kread1_2336 <= tempk1_1_2307 when (read_k_2284_delayed_1_0_2330(0) /=  '0') else tempk2_1_2319;
    -- flow-through select operator MUX_2344_inst
    kread2_2345 <= tempk1_2_2311 when (read_k_2290_delayed_1_0_2339(0) /=  '0') else tempk2_2_2323;
    -- flow-through select operator MUX_2353_inst
    kread3_2354 <= tempk1_3_2315 when (read_k_2296_delayed_1_0_2348(0) /=  '0') else tempk2_3_2327;
    -- flow-through select operator MUX_3031_inst
    n_chl_3032 <= konst_3027_wire_constant when (chl_done_2965(0) /=  '0') else ADD_u16_u16_3030_wire;
    -- flow-through select operator MUX_3040_inst
    MUX_3040_wire <= konst_3036_wire_constant when (num_done_2972(0) /=  '0') else ADD_u2_u2_3039_wire;
    -- flow-through select operator MUX_3042_inst
    n_num_3043 <= MUX_3040_wire when (chl_done_2965(0) /=  '0') else num_1913;
    -- flow-through select operator MUX_3051_inst
    MUX_3051_wire <= konst_3047_wire_constant when (col_done_2977(0) /=  '0') else ADD_u16_u16_3050_wire;
    -- flow-through select operator MUX_3053_inst
    n_col_3054 <= MUX_3051_wire when (num_done_2972(0) /=  '0') else col_1908;
    -- flow-through select operator MUX_3061_inst
    n_row_3062 <= ADD_u16_u16_3059_wire when (row_done_2982(0) /=  '0') else row_1903;
    -- flow-through select operator MUX_3070_inst
    nacc1_3071 <= konst_3068_wire_constant when (num_done_2992_delayed_2_0_3065(0) /=  '0') else acc_val1_2948;
    -- flow-through select operator MUX_3079_inst
    nacc2_3080 <= konst_3077_wire_constant when (num_done_2998_delayed_2_0_3074(0) /=  '0') else acc_val2_2960;
    slice_2041_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2041_inst_req_0;
      slice_2041_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2041_inst_req_1;
      slice_2041_inst_ack_1<= update_ack(0);
      slice_2041_inst: SliceSplitProtocol generic map(name => "slice_2041_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir1_1_2042, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2045_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2045_inst_req_0;
      slice_2045_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2045_inst_req_1;
      slice_2045_inst_ack_1<= update_ack(0);
      slice_2045_inst: SliceSplitProtocol generic map(name => "slice_2045_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir2_1_2046, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2049_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2049_inst_req_0;
      slice_2049_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2049_inst_req_1;
      slice_2049_inst_ack_1<= update_ack(0);
      slice_2049_inst: SliceSplitProtocol generic map(name => "slice_2049_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir3_1_2050, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2053_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2053_inst_req_0;
      slice_2053_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2053_inst_req_1;
      slice_2053_inst_ack_1<= update_ack(0);
      slice_2053_inst: SliceSplitProtocol generic map(name => "slice_2053_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir4_1_2054, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2057_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2057_inst_req_0;
      slice_2057_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2057_inst_req_1;
      slice_2057_inst_ack_1<= update_ack(0);
      slice_2057_inst: SliceSplitProtocol generic map(name => "slice_2057_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir5_1_2058, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2061_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2061_inst_req_0;
      slice_2061_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2061_inst_req_1;
      slice_2061_inst_ack_1<= update_ack(0);
      slice_2061_inst: SliceSplitProtocol generic map(name => "slice_2061_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir6_1_2062, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2065_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2065_inst_req_0;
      slice_2065_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2065_inst_req_1;
      slice_2065_inst_ack_1<= update_ack(0);
      slice_2065_inst: SliceSplitProtocol generic map(name => "slice_2065_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir7_1_2066, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2069_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2069_inst_req_0;
      slice_2069_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2069_inst_req_1;
      slice_2069_inst_ack_1<= update_ack(0);
      slice_2069_inst: SliceSplitProtocol generic map(name => "slice_2069_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread1_1974, dout => ir8_1_2070, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2073_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2073_inst_req_0;
      slice_2073_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2073_inst_req_1;
      slice_2073_inst_ack_1<= update_ack(0);
      slice_2073_inst: SliceSplitProtocol generic map(name => "slice_2073_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir1_2_2074, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2077_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2077_inst_req_0;
      slice_2077_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2077_inst_req_1;
      slice_2077_inst_ack_1<= update_ack(0);
      slice_2077_inst: SliceSplitProtocol generic map(name => "slice_2077_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir2_2_2078, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2081_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2081_inst_req_0;
      slice_2081_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2081_inst_req_1;
      slice_2081_inst_ack_1<= update_ack(0);
      slice_2081_inst: SliceSplitProtocol generic map(name => "slice_2081_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir3_2_2082, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2085_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2085_inst_req_0;
      slice_2085_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2085_inst_req_1;
      slice_2085_inst_ack_1<= update_ack(0);
      slice_2085_inst: SliceSplitProtocol generic map(name => "slice_2085_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir4_2_2086, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2089_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2089_inst_req_0;
      slice_2089_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2089_inst_req_1;
      slice_2089_inst_ack_1<= update_ack(0);
      slice_2089_inst: SliceSplitProtocol generic map(name => "slice_2089_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir5_2_2090, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2093_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2093_inst_req_0;
      slice_2093_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2093_inst_req_1;
      slice_2093_inst_ack_1<= update_ack(0);
      slice_2093_inst: SliceSplitProtocol generic map(name => "slice_2093_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir6_2_2094, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2097_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2097_inst_req_0;
      slice_2097_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2097_inst_req_1;
      slice_2097_inst_ack_1<= update_ack(0);
      slice_2097_inst: SliceSplitProtocol generic map(name => "slice_2097_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir7_2_2098, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2101_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2101_inst_req_0;
      slice_2101_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2101_inst_req_1;
      slice_2101_inst_ack_1<= update_ack(0);
      slice_2101_inst: SliceSplitProtocol generic map(name => "slice_2101_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread2_1983, dout => ir8_2_2102, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2105_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2105_inst_req_0;
      slice_2105_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2105_inst_req_1;
      slice_2105_inst_ack_1<= update_ack(0);
      slice_2105_inst: SliceSplitProtocol generic map(name => "slice_2105_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir1_3_2106, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2109_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2109_inst_req_0;
      slice_2109_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2109_inst_req_1;
      slice_2109_inst_ack_1<= update_ack(0);
      slice_2109_inst: SliceSplitProtocol generic map(name => "slice_2109_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir2_3_2110, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2113_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2113_inst_req_0;
      slice_2113_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2113_inst_req_1;
      slice_2113_inst_ack_1<= update_ack(0);
      slice_2113_inst: SliceSplitProtocol generic map(name => "slice_2113_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir3_3_2114, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2117_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2117_inst_req_0;
      slice_2117_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2117_inst_req_1;
      slice_2117_inst_ack_1<= update_ack(0);
      slice_2117_inst: SliceSplitProtocol generic map(name => "slice_2117_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir4_3_2118, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2121_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2121_inst_req_0;
      slice_2121_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2121_inst_req_1;
      slice_2121_inst_ack_1<= update_ack(0);
      slice_2121_inst: SliceSplitProtocol generic map(name => "slice_2121_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir5_3_2122, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2125_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2125_inst_req_0;
      slice_2125_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2125_inst_req_1;
      slice_2125_inst_ack_1<= update_ack(0);
      slice_2125_inst: SliceSplitProtocol generic map(name => "slice_2125_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir6_3_2126, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2129_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2129_inst_req_0;
      slice_2129_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2129_inst_req_1;
      slice_2129_inst_ack_1<= update_ack(0);
      slice_2129_inst: SliceSplitProtocol generic map(name => "slice_2129_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir7_3_2130, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2133_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2133_inst_req_0;
      slice_2133_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2133_inst_req_1;
      slice_2133_inst_ack_1<= update_ack(0);
      slice_2133_inst: SliceSplitProtocol generic map(name => "slice_2133_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread3_1992, dout => ir8_3_2134, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2137_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2137_inst_req_0;
      slice_2137_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2137_inst_req_1;
      slice_2137_inst_ack_1<= update_ack(0);
      slice_2137_inst: SliceSplitProtocol generic map(name => "slice_2137_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir1_4_2138, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2141_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2141_inst_req_0;
      slice_2141_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2141_inst_req_1;
      slice_2141_inst_ack_1<= update_ack(0);
      slice_2141_inst: SliceSplitProtocol generic map(name => "slice_2141_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir2_4_2142, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2145_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2145_inst_req_0;
      slice_2145_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2145_inst_req_1;
      slice_2145_inst_ack_1<= update_ack(0);
      slice_2145_inst: SliceSplitProtocol generic map(name => "slice_2145_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir3_4_2146, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2149_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2149_inst_req_0;
      slice_2149_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2149_inst_req_1;
      slice_2149_inst_ack_1<= update_ack(0);
      slice_2149_inst: SliceSplitProtocol generic map(name => "slice_2149_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir4_4_2150, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2153_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2153_inst_req_0;
      slice_2153_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2153_inst_req_1;
      slice_2153_inst_ack_1<= update_ack(0);
      slice_2153_inst: SliceSplitProtocol generic map(name => "slice_2153_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir5_4_2154, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2157_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2157_inst_req_0;
      slice_2157_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2157_inst_req_1;
      slice_2157_inst_ack_1<= update_ack(0);
      slice_2157_inst: SliceSplitProtocol generic map(name => "slice_2157_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir6_4_2158, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2161_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2161_inst_req_0;
      slice_2161_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2161_inst_req_1;
      slice_2161_inst_ack_1<= update_ack(0);
      slice_2161_inst: SliceSplitProtocol generic map(name => "slice_2161_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir7_4_2162, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2165_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2165_inst_req_0;
      slice_2165_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2165_inst_req_1;
      slice_2165_inst_ack_1<= update_ack(0);
      slice_2165_inst: SliceSplitProtocol generic map(name => "slice_2165_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => iread4_2001, dout => ir8_4_2166, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2357_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2357_inst_req_0;
      slice_2357_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2357_inst_req_1;
      slice_2357_inst_ack_1<= update_ack(0);
      slice_2357_inst: SliceSplitProtocol generic map(name => "slice_2357_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr1_1_2358, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2361_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2361_inst_req_0;
      slice_2361_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2361_inst_req_1;
      slice_2361_inst_ack_1<= update_ack(0);
      slice_2361_inst: SliceSplitProtocol generic map(name => "slice_2361_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr2_1_2362, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2365_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2365_inst_req_0;
      slice_2365_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2365_inst_req_1;
      slice_2365_inst_ack_1<= update_ack(0);
      slice_2365_inst: SliceSplitProtocol generic map(name => "slice_2365_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr3_1_2366, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2369_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2369_inst_req_0;
      slice_2369_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2369_inst_req_1;
      slice_2369_inst_ack_1<= update_ack(0);
      slice_2369_inst: SliceSplitProtocol generic map(name => "slice_2369_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr4_1_2370, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2373_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2373_inst_req_0;
      slice_2373_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2373_inst_req_1;
      slice_2373_inst_ack_1<= update_ack(0);
      slice_2373_inst: SliceSplitProtocol generic map(name => "slice_2373_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr5_1_2374, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2377_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2377_inst_req_0;
      slice_2377_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2377_inst_req_1;
      slice_2377_inst_ack_1<= update_ack(0);
      slice_2377_inst: SliceSplitProtocol generic map(name => "slice_2377_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr6_1_2378, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2381_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2381_inst_req_0;
      slice_2381_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2381_inst_req_1;
      slice_2381_inst_ack_1<= update_ack(0);
      slice_2381_inst: SliceSplitProtocol generic map(name => "slice_2381_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr7_1_2382, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2385_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2385_inst_req_0;
      slice_2385_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2385_inst_req_1;
      slice_2385_inst_ack_1<= update_ack(0);
      slice_2385_inst: SliceSplitProtocol generic map(name => "slice_2385_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread1_2336, dout => kr8_1_2386, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2389_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2389_inst_req_0;
      slice_2389_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2389_inst_req_1;
      slice_2389_inst_ack_1<= update_ack(0);
      slice_2389_inst: SliceSplitProtocol generic map(name => "slice_2389_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr1_2_2390, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2393_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2393_inst_req_0;
      slice_2393_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2393_inst_req_1;
      slice_2393_inst_ack_1<= update_ack(0);
      slice_2393_inst: SliceSplitProtocol generic map(name => "slice_2393_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr2_2_2394, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2397_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2397_inst_req_0;
      slice_2397_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2397_inst_req_1;
      slice_2397_inst_ack_1<= update_ack(0);
      slice_2397_inst: SliceSplitProtocol generic map(name => "slice_2397_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr3_2_2398, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2401_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2401_inst_req_0;
      slice_2401_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2401_inst_req_1;
      slice_2401_inst_ack_1<= update_ack(0);
      slice_2401_inst: SliceSplitProtocol generic map(name => "slice_2401_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr4_2_2402, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2405_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2405_inst_req_0;
      slice_2405_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2405_inst_req_1;
      slice_2405_inst_ack_1<= update_ack(0);
      slice_2405_inst: SliceSplitProtocol generic map(name => "slice_2405_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr5_2_2406, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2409_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2409_inst_req_0;
      slice_2409_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2409_inst_req_1;
      slice_2409_inst_ack_1<= update_ack(0);
      slice_2409_inst: SliceSplitProtocol generic map(name => "slice_2409_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr6_2_2410, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2413_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2413_inst_req_0;
      slice_2413_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2413_inst_req_1;
      slice_2413_inst_ack_1<= update_ack(0);
      slice_2413_inst: SliceSplitProtocol generic map(name => "slice_2413_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr7_2_2414, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2417_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2417_inst_req_0;
      slice_2417_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2417_inst_req_1;
      slice_2417_inst_ack_1<= update_ack(0);
      slice_2417_inst: SliceSplitProtocol generic map(name => "slice_2417_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread2_2345, dout => kr8_2_2418, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2421_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2421_inst_req_0;
      slice_2421_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2421_inst_req_1;
      slice_2421_inst_ack_1<= update_ack(0);
      slice_2421_inst: SliceSplitProtocol generic map(name => "slice_2421_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr1_3_2422, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2425_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2425_inst_req_0;
      slice_2425_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2425_inst_req_1;
      slice_2425_inst_ack_1<= update_ack(0);
      slice_2425_inst: SliceSplitProtocol generic map(name => "slice_2425_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr2_3_2426, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2429_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2429_inst_req_0;
      slice_2429_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2429_inst_req_1;
      slice_2429_inst_ack_1<= update_ack(0);
      slice_2429_inst: SliceSplitProtocol generic map(name => "slice_2429_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr3_3_2430, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2433_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2433_inst_req_0;
      slice_2433_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2433_inst_req_1;
      slice_2433_inst_ack_1<= update_ack(0);
      slice_2433_inst: SliceSplitProtocol generic map(name => "slice_2433_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr4_3_2434, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2437_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2437_inst_req_0;
      slice_2437_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2437_inst_req_1;
      slice_2437_inst_ack_1<= update_ack(0);
      slice_2437_inst: SliceSplitProtocol generic map(name => "slice_2437_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr5_3_2438, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2441_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2441_inst_req_0;
      slice_2441_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2441_inst_req_1;
      slice_2441_inst_ack_1<= update_ack(0);
      slice_2441_inst: SliceSplitProtocol generic map(name => "slice_2441_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr6_3_2442, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2445_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2445_inst_req_0;
      slice_2445_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2445_inst_req_1;
      slice_2445_inst_ack_1<= update_ack(0);
      slice_2445_inst: SliceSplitProtocol generic map(name => "slice_2445_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr7_3_2446, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_2449_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_2449_inst_req_0;
      slice_2449_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_2449_inst_req_1;
      slice_2449_inst_ack_1<= update_ack(0);
      slice_2449_inst: SliceSplitProtocol generic map(name => "slice_2449_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 2, flow_through => false,  full_rate => true) -- 
        port map( din => kread3_2354, dout => kr8_3_2450, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_acc1_2884_delayed_2_0_2937_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc1_2884_delayed_2_0_2937_inst_req_0;
      W_acc1_2884_delayed_2_0_2937_inst_ack_0<= wack(0);
      rreq(0) <= W_acc1_2884_delayed_2_0_2937_inst_req_1;
      W_acc1_2884_delayed_2_0_2937_inst_ack_1<= rack(0);
      W_acc1_2884_delayed_2_0_2937_inst : InterlockBuffer generic map ( -- 
        name => "W_acc1_2884_delayed_2_0_2937_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc1_1892,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc1_2884_delayed_2_0_2939,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_acc2_2893_delayed_2_0_2949_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_acc2_2893_delayed_2_0_2949_inst_req_0;
      W_acc2_2893_delayed_2_0_2949_inst_ack_0<= wack(0);
      rreq(0) <= W_acc2_2893_delayed_2_0_2949_inst_req_1;
      W_acc2_2893_delayed_2_0_2949_inst_ack_1<= rack(0);
      W_acc2_2893_delayed_2_0_2949_inst : InterlockBuffer generic map ( -- 
        name => "W_acc2_2893_delayed_2_0_2949_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => acc2_1898,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => acc2_2893_delayed_2_0_2951,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2992_delayed_2_0_3063_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2992_delayed_2_0_3063_inst_req_0;
      W_num_done_2992_delayed_2_0_3063_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2992_delayed_2_0_3063_inst_req_1;
      W_num_done_2992_delayed_2_0_3063_inst_ack_1<= rack(0);
      W_num_done_2992_delayed_2_0_3063_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2992_delayed_2_0_3063_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2992_delayed_2_0_3065,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_2998_delayed_2_0_3072_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_2998_delayed_2_0_3072_inst_req_0;
      W_num_done_2998_delayed_2_0_3072_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_2998_delayed_2_0_3072_inst_req_1;
      W_num_done_2998_delayed_2_0_3072_inst_ack_1<= rack(0);
      W_num_done_2998_delayed_2_0_3072_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_2998_delayed_2_0_3072_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_2998_delayed_2_0_3074,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_num_done_3003_delayed_2_0_3081_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_num_done_3003_delayed_2_0_3081_inst_req_0;
      W_num_done_3003_delayed_2_0_3081_inst_ack_0<= wack(0);
      rreq(0) <= W_num_done_3003_delayed_2_0_3081_inst_req_1;
      W_num_done_3003_delayed_2_0_3081_inst_ack_1<= rack(0);
      W_num_done_3003_delayed_2_0_3081_inst : InterlockBuffer generic map ( -- 
        name => "W_num_done_3003_delayed_2_0_3081_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => num_done_2972,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => num_done_3003_delayed_2_0_3083,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1946_delayed_1_0_1966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1946_delayed_1_0_1966_inst_req_0;
      W_read_ip_1946_delayed_1_0_1966_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1946_delayed_1_0_1966_inst_req_1;
      W_read_ip_1946_delayed_1_0_1966_inst_ack_1<= rack(0);
      W_read_ip_1946_delayed_1_0_1966_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1946_delayed_1_0_1966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1946_delayed_1_0_1968,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1952_delayed_1_0_1975_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1952_delayed_1_0_1975_inst_req_0;
      W_read_ip_1952_delayed_1_0_1975_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1952_delayed_1_0_1975_inst_req_1;
      W_read_ip_1952_delayed_1_0_1975_inst_ack_1<= rack(0);
      W_read_ip_1952_delayed_1_0_1975_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1952_delayed_1_0_1975_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1952_delayed_1_0_1977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1958_delayed_1_0_1984_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1958_delayed_1_0_1984_inst_req_0;
      W_read_ip_1958_delayed_1_0_1984_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1958_delayed_1_0_1984_inst_req_1;
      W_read_ip_1958_delayed_1_0_1984_inst_ack_1<= rack(0);
      W_read_ip_1958_delayed_1_0_1984_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1958_delayed_1_0_1984_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1958_delayed_1_0_1986,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_ip_1964_delayed_1_0_1993_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_ip_1964_delayed_1_0_1993_inst_req_0;
      W_read_ip_1964_delayed_1_0_1993_inst_ack_0<= wack(0);
      rreq(0) <= W_read_ip_1964_delayed_1_0_1993_inst_req_1;
      W_read_ip_1964_delayed_1_0_1993_inst_ack_1<= rack(0);
      W_read_ip_1964_delayed_1_0_1993_inst : InterlockBuffer generic map ( -- 
        name => "W_read_ip_1964_delayed_1_0_1993_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_ip_1933,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_ip_1964_delayed_1_0_1995,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2284_delayed_1_0_2328_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2284_delayed_1_0_2328_inst_req_0;
      W_read_k_2284_delayed_1_0_2328_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2284_delayed_1_0_2328_inst_req_1;
      W_read_k_2284_delayed_1_0_2328_inst_ack_1<= rack(0);
      W_read_k_2284_delayed_1_0_2328_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2284_delayed_1_0_2328_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2284_delayed_1_0_2330,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2290_delayed_1_0_2337_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2290_delayed_1_0_2337_inst_req_0;
      W_read_k_2290_delayed_1_0_2337_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2290_delayed_1_0_2337_inst_req_1;
      W_read_k_2290_delayed_1_0_2337_inst_ack_1<= rack(0);
      W_read_k_2290_delayed_1_0_2337_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2290_delayed_1_0_2337_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2290_delayed_1_0_2339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_read_k_2296_delayed_1_0_2346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_k_2296_delayed_1_0_2346_inst_req_0;
      W_read_k_2296_delayed_1_0_2346_inst_ack_0<= wack(0);
      rreq(0) <= W_read_k_2296_delayed_1_0_2346_inst_req_1;
      W_read_k_2296_delayed_1_0_2346_inst_ack_1<= rack(0);
      W_read_k_2296_delayed_1_0_2346_inst : InterlockBuffer generic map ( -- 
        name => "W_read_k_2296_delayed_1_0_2346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_k_2303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_k_2296_delayed_1_0_2348,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2941_delayed_1_0_3004_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2941_delayed_1_0_3004_inst_req_0;
      W_store_kernel_2941_delayed_1_0_3004_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2941_delayed_1_0_3004_inst_req_1;
      W_store_kernel_2941_delayed_1_0_3004_inst_ack_1<= rack(0);
      W_store_kernel_2941_delayed_1_0_3004_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2941_delayed_1_0_3004_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2941_delayed_1_0_3006,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2945_delayed_1_0_3011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2945_delayed_1_0_3011_inst_req_0;
      W_store_kernel_2945_delayed_1_0_3011_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2945_delayed_1_0_3011_inst_req_1;
      W_store_kernel_2945_delayed_1_0_3011_inst_ack_1<= rack(0);
      W_store_kernel_2945_delayed_1_0_3011_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2945_delayed_1_0_3011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2945_delayed_1_0_3013,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_store_kernel_2949_delayed_1_0_3018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_store_kernel_2949_delayed_1_0_3018_inst_req_0;
      W_store_kernel_2949_delayed_1_0_3018_inst_ack_0<= wack(0);
      rreq(0) <= W_store_kernel_2949_delayed_1_0_3018_inst_req_1;
      W_store_kernel_2949_delayed_1_0_3018_inst_ack_1<= rack(0);
      W_store_kernel_2949_delayed_1_0_3018_inst : InterlockBuffer generic map ( -- 
        name => "W_store_kernel_2949_delayed_1_0_3018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => store_kernel_2998,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => store_kernel_2949_delayed_1_0_3020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1978_delayed_1_0_2011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1978_delayed_1_0_2011_inst_req_0;
      W_write_input_1978_delayed_1_0_2011_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1978_delayed_1_0_2011_inst_req_1;
      W_write_input_1978_delayed_1_0_2011_inst_ack_1<= rack(0);
      W_write_input_1978_delayed_1_0_2011_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1978_delayed_1_0_2011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1978_delayed_1_0_2013,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1982_delayed_1_0_2018_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1982_delayed_1_0_2018_inst_req_0;
      W_write_input_1982_delayed_1_0_2018_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1982_delayed_1_0_2018_inst_req_1;
      W_write_input_1982_delayed_1_0_2018_inst_ack_1<= rack(0);
      W_write_input_1982_delayed_1_0_2018_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1982_delayed_1_0_2018_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1982_delayed_1_0_2020,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1986_delayed_1_0_2025_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1986_delayed_1_0_2025_inst_req_0;
      W_write_input_1986_delayed_1_0_2025_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1986_delayed_1_0_2025_inst_req_1;
      W_write_input_1986_delayed_1_0_2025_inst_ack_1<= rack(0);
      W_write_input_1986_delayed_1_0_2025_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1986_delayed_1_0_2025_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1986_delayed_1_0_2027,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_input_1990_delayed_1_0_2032_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_input_1990_delayed_1_0_2032_inst_req_0;
      W_write_input_1990_delayed_1_0_2032_inst_ack_0<= wack(0);
      rreq(0) <= W_write_input_1990_delayed_1_0_2032_inst_req_1;
      W_write_input_1990_delayed_1_0_2032_inst_ack_1<= rack(0);
      W_write_input_1990_delayed_1_0_2032_inst : InterlockBuffer generic map ( -- 
        name => "W_write_input_1990_delayed_1_0_2032_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_input_2010,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_input_1990_delayed_1_0_2034,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3032_1923_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3032_1923_buf_req_0;
      n_chl_3032_1923_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3032_1923_buf_req_1;
      n_chl_3032_1923_buf_ack_1<= rack(0);
      n_chl_3032_1923_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3032_1923_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3032,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3032_1923_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3054_1912_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3054_1912_buf_req_0;
      n_col_3054_1912_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3054_1912_buf_req_1;
      n_col_3054_1912_buf_ack_1<= rack(0);
      n_col_3054_1912_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3054_1912_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3054,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3054_1912_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_num_3043_1918_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_num_3043_1918_buf_req_0;
      n_num_3043_1918_buf_ack_0<= wack(0);
      rreq(0) <= n_num_3043_1918_buf_req_1;
      n_num_3043_1918_buf_ack_1<= rack(0);
      n_num_3043_1918_buf : InterlockBuffer generic map ( -- 
        name => "n_num_3043_1918_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_num_3043,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_num_3043_1918_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3062_1907_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3062_1907_buf_req_0;
      n_row_3062_1907_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3062_1907_buf_req_1;
      n_row_3062_1907_buf_ack_1<= rack(0);
      n_row_3062_1907_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3062_1907_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3062,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3062_1907_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc1_3071_1897_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc1_3071_1897_buf_req_0;
      nacc1_3071_1897_buf_ack_0<= wack(0);
      rreq(0) <= nacc1_3071_1897_buf_req_1;
      nacc1_3071_1897_buf_ack_1<= rack(0);
      nacc1_3071_1897_buf : InterlockBuffer generic map ( -- 
        name => "nacc1_3071_1897_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc1_3071,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc1_3071_1897_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nacc2_3080_1902_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nacc2_3080_1902_buf_req_0;
      nacc2_3080_1902_buf_ack_0<= wack(0);
      rreq(0) <= nacc2_3080_1902_buf_req_1;
      nacc2_3080_1902_buf_ack_1<= rack(0);
      nacc2_3080_1902_buf : InterlockBuffer generic map ( -- 
        name => "nacc2_3080_1902_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nacc2_3080,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nacc2_3080_1902_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2169_inst
    process(ir1_1_2042) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir1_1_2042(7 downto 0);
      ival1_1_2170 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2173_inst
    process(ir2_1_2046) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir2_1_2046(7 downto 0);
      ival2_1_2174 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2177_inst
    process(ir3_1_2050) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir3_1_2050(7 downto 0);
      ival3_1_2178 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2181_inst
    process(ir4_1_2054) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir4_1_2054(7 downto 0);
      ival4_1_2182 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2185_inst
    process(ir5_1_2058) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir5_1_2058(7 downto 0);
      ival5_1_2186 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2189_inst
    process(ir6_1_2062) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir6_1_2062(7 downto 0);
      ival6_1_2190 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2193_inst
    process(ir7_1_2066) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir7_1_2066(7 downto 0);
      ival7_1_2194 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2197_inst
    process(ir8_1_2070) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir8_1_2070(7 downto 0);
      ival8_1_2198 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2201_inst
    process(ir1_2_2074) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir1_2_2074(7 downto 0);
      ival1_2_2202 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2205_inst
    process(ir2_2_2078) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir2_2_2078(7 downto 0);
      ival2_2_2206 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2209_inst
    process(ir3_2_2082) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir3_2_2082(7 downto 0);
      ival3_2_2210 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2213_inst
    process(ir4_2_2086) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir4_2_2086(7 downto 0);
      ival4_2_2214 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2217_inst
    process(ir5_2_2090) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir5_2_2090(7 downto 0);
      ival5_2_2218 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2221_inst
    process(ir6_2_2094) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir6_2_2094(7 downto 0);
      ival6_2_2222 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2225_inst
    process(ir7_2_2098) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir7_2_2098(7 downto 0);
      ival7_2_2226 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2229_inst
    process(ir8_2_2102) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir8_2_2102(7 downto 0);
      ival8_2_2230 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2233_inst
    process(ir1_3_2106) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir1_3_2106(7 downto 0);
      ival1_3_2234 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2237_inst
    process(ir2_3_2110) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir2_3_2110(7 downto 0);
      ival2_3_2238 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2241_inst
    process(ir3_3_2114) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir3_3_2114(7 downto 0);
      ival3_3_2242 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2245_inst
    process(ir4_3_2118) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir4_3_2118(7 downto 0);
      ival4_3_2246 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2249_inst
    process(ir5_3_2122) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir5_3_2122(7 downto 0);
      ival5_3_2250 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2253_inst
    process(ir6_3_2126) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir6_3_2126(7 downto 0);
      ival6_3_2254 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2257_inst
    process(ir7_3_2130) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir7_3_2130(7 downto 0);
      ival7_3_2258 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2261_inst
    process(ir8_3_2134) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir8_3_2134(7 downto 0);
      ival8_3_2262 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2265_inst
    process(ir1_4_2138) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir1_4_2138(7 downto 0);
      ival1_4_2266 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2269_inst
    process(ir2_4_2142) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir2_4_2142(7 downto 0);
      ival2_4_2270 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2273_inst
    process(ir3_4_2146) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir3_4_2146(7 downto 0);
      ival3_4_2274 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2277_inst
    process(ir4_4_2150) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir4_4_2150(7 downto 0);
      ival4_4_2278 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2281_inst
    process(ir5_4_2154) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir5_4_2154(7 downto 0);
      ival5_4_2282 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2285_inst
    process(ir6_4_2158) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir6_4_2158(7 downto 0);
      ival6_4_2286 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2289_inst
    process(ir7_4_2162) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir7_4_2162(7 downto 0);
      ival7_4_2290 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2293_inst
    process(ir8_4_2166) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ir8_4_2166(7 downto 0);
      ival8_4_2294 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2453_inst
    process(kr1_1_2358) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr1_1_2358(7 downto 0);
      kval1_1_2454 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2457_inst
    process(kr2_1_2362) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr2_1_2362(7 downto 0);
      kval2_1_2458 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2461_inst
    process(kr3_1_2366) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr3_1_2366(7 downto 0);
      kval3_1_2462 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2465_inst
    process(kr4_1_2370) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr4_1_2370(7 downto 0);
      kval4_1_2466 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2469_inst
    process(kr5_1_2374) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr5_1_2374(7 downto 0);
      kval5_1_2470 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2473_inst
    process(kr6_1_2378) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr6_1_2378(7 downto 0);
      kval6_1_2474 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2477_inst
    process(kr7_1_2382) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr7_1_2382(7 downto 0);
      kval7_1_2478 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2481_inst
    process(kr8_1_2386) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr8_1_2386(7 downto 0);
      kval8_1_2482 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2485_inst
    process(kr1_2_2390) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr1_2_2390(7 downto 0);
      kval1_2_2486 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2489_inst
    process(kr2_2_2394) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr2_2_2394(7 downto 0);
      kval2_2_2490 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2493_inst
    process(kr3_2_2398) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr3_2_2398(7 downto 0);
      kval3_2_2494 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2497_inst
    process(kr4_2_2402) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr4_2_2402(7 downto 0);
      kval4_2_2498 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2501_inst
    process(kr5_2_2406) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr5_2_2406(7 downto 0);
      kval5_2_2502 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2505_inst
    process(kr6_2_2410) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr6_2_2410(7 downto 0);
      kval6_2_2506 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2509_inst
    process(kr7_2_2414) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr7_2_2414(7 downto 0);
      kval7_2_2510 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2513_inst
    process(kr8_2_2418) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr8_2_2418(7 downto 0);
      kval8_2_2514 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2517_inst
    process(kr1_3_2422) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr1_3_2422(7 downto 0);
      kval1_3_2518 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2521_inst
    process(kr2_3_2426) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr2_3_2426(7 downto 0);
      kval2_3_2522 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2525_inst
    process(kr3_3_2430) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr3_3_2430(7 downto 0);
      kval3_3_2526 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2529_inst
    process(kr4_3_2434) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr4_3_2434(7 downto 0);
      kval4_3_2530 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2533_inst
    process(kr5_3_2438) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr5_3_2438(7 downto 0);
      kval5_3_2534 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2537_inst
    process(kr6_3_2442) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr6_3_2442(7 downto 0);
      kval6_3_2538 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2541_inst
    process(kr7_3_2446) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr7_3_2446(7 downto 0);
      kval7_3_2542 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2545_inst
    process(kr8_3_2450) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := kr8_3_2450(7 downto 0);
      kval8_3_2546 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2551_inst
    process(MUL_i8_i8_2550_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2550_wire(7 downto 0);
      mul_val1_1_2552 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2557_inst
    process(MUL_i8_i8_2556_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2556_wire(7 downto 0);
      mul_val2_1_2558 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2563_inst
    process(MUL_i8_i8_2562_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2562_wire(7 downto 0);
      mul_val3_1_2564 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2569_inst
    process(MUL_i8_i8_2568_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2568_wire(7 downto 0);
      mul_val4_1_2570 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2575_inst
    process(MUL_i8_i8_2574_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2574_wire(7 downto 0);
      mul_val5_1_2576 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2581_inst
    process(MUL_i8_i8_2580_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2580_wire(7 downto 0);
      mul_val6_1_2582 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2587_inst
    process(MUL_i8_i8_2586_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2586_wire(7 downto 0);
      mul_val7_1_2588 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2593_inst
    process(MUL_i8_i8_2592_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2592_wire(7 downto 0);
      mul_val8_1_2594 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2599_inst
    process(MUL_i8_i8_2598_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2598_wire(7 downto 0);
      mul_val1_2_2600 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2605_inst
    process(MUL_i8_i8_2604_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2604_wire(7 downto 0);
      mul_val2_2_2606 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2611_inst
    process(MUL_i8_i8_2610_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2610_wire(7 downto 0);
      mul_val3_2_2612 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2617_inst
    process(MUL_i8_i8_2616_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2616_wire(7 downto 0);
      mul_val4_2_2618 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2623_inst
    process(MUL_i8_i8_2622_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2622_wire(7 downto 0);
      mul_val5_2_2624 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2629_inst
    process(MUL_i8_i8_2628_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2628_wire(7 downto 0);
      mul_val6_2_2630 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2635_inst
    process(MUL_i8_i8_2634_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2634_wire(7 downto 0);
      mul_val7_2_2636 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2641_inst
    process(MUL_i8_i8_2640_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2640_wire(7 downto 0);
      mul_val8_2_2642 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2647_inst
    process(MUL_i8_i8_2646_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2646_wire(7 downto 0);
      mul_val1_3_2648 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2653_inst
    process(MUL_i8_i8_2652_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2652_wire(7 downto 0);
      mul_val2_3_2654 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2659_inst
    process(MUL_i8_i8_2658_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2658_wire(7 downto 0);
      mul_val3_3_2660 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2665_inst
    process(MUL_i8_i8_2664_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2664_wire(7 downto 0);
      mul_val4_3_2666 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2671_inst
    process(MUL_i8_i8_2670_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2670_wire(7 downto 0);
      mul_val5_3_2672 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2677_inst
    process(MUL_i8_i8_2676_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2676_wire(7 downto 0);
      mul_val6_3_2678 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2683_inst
    process(MUL_i8_i8_2682_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2682_wire(7 downto 0);
      mul_val7_3_2684 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2689_inst
    process(MUL_i8_i8_2688_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2688_wire(7 downto 0);
      mul_val8_3_2690 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2695_inst
    process(MUL_i8_i8_2694_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2694_wire(7 downto 0);
      mul_val1_4_2696 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2701_inst
    process(MUL_i8_i8_2700_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2700_wire(7 downto 0);
      mul_val2_4_2702 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2707_inst
    process(MUL_i8_i8_2706_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2706_wire(7 downto 0);
      mul_val3_4_2708 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2713_inst
    process(MUL_i8_i8_2712_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2712_wire(7 downto 0);
      mul_val4_4_2714 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2719_inst
    process(MUL_i8_i8_2718_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2718_wire(7 downto 0);
      mul_val5_4_2720 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2725_inst
    process(MUL_i8_i8_2724_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2724_wire(7 downto 0);
      mul_val6_4_2726 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2731_inst
    process(MUL_i8_i8_2730_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2730_wire(7 downto 0);
      mul_val7_4_2732 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2737_inst
    process(MUL_i8_i8_2736_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2736_wire(7 downto 0);
      mul_val8_4_2738 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2743_inst
    process(MUL_i8_i8_2742_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2742_wire(7 downto 0);
      mul_val1_5_2744 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2749_inst
    process(MUL_i8_i8_2748_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2748_wire(7 downto 0);
      mul_val2_5_2750 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2755_inst
    process(MUL_i8_i8_2754_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2754_wire(7 downto 0);
      mul_val3_5_2756 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2761_inst
    process(MUL_i8_i8_2760_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2760_wire(7 downto 0);
      mul_val4_5_2762 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2767_inst
    process(MUL_i8_i8_2766_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2766_wire(7 downto 0);
      mul_val5_5_2768 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2773_inst
    process(MUL_i8_i8_2772_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2772_wire(7 downto 0);
      mul_val6_5_2774 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2779_inst
    process(MUL_i8_i8_2778_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2778_wire(7 downto 0);
      mul_val7_5_2780 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2785_inst
    process(MUL_i8_i8_2784_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2784_wire(7 downto 0);
      mul_val8_5_2786 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2791_inst
    process(MUL_i8_i8_2790_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2790_wire(7 downto 0);
      mul_val1_6_2792 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2797_inst
    process(MUL_i8_i8_2796_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2796_wire(7 downto 0);
      mul_val2_6_2798 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2803_inst
    process(MUL_i8_i8_2802_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2802_wire(7 downto 0);
      mul_val3_6_2804 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2809_inst
    process(MUL_i8_i8_2808_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2808_wire(7 downto 0);
      mul_val4_6_2810 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2815_inst
    process(MUL_i8_i8_2814_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2814_wire(7 downto 0);
      mul_val5_6_2816 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2821_inst
    process(MUL_i8_i8_2820_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2820_wire(7 downto 0);
      mul_val6_6_2822 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2827_inst
    process(MUL_i8_i8_2826_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2826_wire(7 downto 0);
      mul_val7_6_2828 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2833_inst
    process(MUL_i8_i8_2832_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := MUL_i8_i8_2832_wire(7 downto 0);
      mul_val8_6_2834 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3087_inst
    process(acc_val1_2948) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := acc_val1_2948(7 downto 0);
      type_cast_3087_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3089_inst
    process(acc_val2_2960) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := acc_val2_2960(7 downto 0);
      type_cast_3089_wire <= tmp_var; -- 
    end process;
    do_while_stmt_1890_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_3094_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1890_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1890_branch_req_0,
          ack0 => do_while_stmt_1890_branch_ack_0,
          ack1 => do_while_stmt_1890_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_i8_i8_2838_inst
    process(mul_val1_1_2552, mul_val2_1_2558) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_1_2552, mul_val2_1_2558, tmp_var);
      ADD_i8_i8_2838_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2841_inst
    process(mul_val3_1_2564, mul_val4_1_2570) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_1_2564, mul_val4_1_2570, tmp_var);
      ADD_i8_i8_2841_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2842_inst
    process(ADD_i8_i8_2838_wire, ADD_i8_i8_2841_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2838_wire, ADD_i8_i8_2841_wire, tmp_var);
      ADD_i8_i8_2842_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2845_inst
    process(mul_val5_1_2576, mul_val6_1_2582) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_1_2576, mul_val6_1_2582, tmp_var);
      ADD_i8_i8_2845_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2848_inst
    process(mul_val7_1_2588, mul_val8_1_2594) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_1_2588, mul_val8_1_2594, tmp_var);
      ADD_i8_i8_2848_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2849_inst
    process(ADD_i8_i8_2845_wire, ADD_i8_i8_2848_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2845_wire, ADD_i8_i8_2848_wire, tmp_var);
      ADD_i8_i8_2849_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2850_inst
    process(ADD_i8_i8_2842_wire, ADD_i8_i8_2849_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2842_wire, ADD_i8_i8_2849_wire, tmp_var);
      t_acc_val1_2851 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2855_inst
    process(mul_val1_2_2600, mul_val2_2_2606) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_2_2600, mul_val2_2_2606, tmp_var);
      ADD_i8_i8_2855_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2858_inst
    process(mul_val3_2_2612, mul_val4_2_2618) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_2_2612, mul_val4_2_2618, tmp_var);
      ADD_i8_i8_2858_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2859_inst
    process(ADD_i8_i8_2855_wire, ADD_i8_i8_2858_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2855_wire, ADD_i8_i8_2858_wire, tmp_var);
      ADD_i8_i8_2859_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2862_inst
    process(mul_val5_2_2624, mul_val6_2_2630) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_2_2624, mul_val6_2_2630, tmp_var);
      ADD_i8_i8_2862_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2865_inst
    process(mul_val7_2_2636, mul_val8_2_2642) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_2_2636, mul_val8_2_2642, tmp_var);
      ADD_i8_i8_2865_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2866_inst
    process(ADD_i8_i8_2862_wire, ADD_i8_i8_2865_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2862_wire, ADD_i8_i8_2865_wire, tmp_var);
      ADD_i8_i8_2866_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2867_inst
    process(ADD_i8_i8_2859_wire, ADD_i8_i8_2866_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2859_wire, ADD_i8_i8_2866_wire, tmp_var);
      t_acc_val2_2868 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2872_inst
    process(mul_val1_3_2648, mul_val2_3_2654) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_3_2648, mul_val2_3_2654, tmp_var);
      ADD_i8_i8_2872_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2875_inst
    process(mul_val3_3_2660, mul_val4_3_2666) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_3_2660, mul_val4_3_2666, tmp_var);
      ADD_i8_i8_2875_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2876_inst
    process(ADD_i8_i8_2872_wire, ADD_i8_i8_2875_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2872_wire, ADD_i8_i8_2875_wire, tmp_var);
      ADD_i8_i8_2876_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2879_inst
    process(mul_val5_3_2672, mul_val6_3_2678) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_3_2672, mul_val6_3_2678, tmp_var);
      ADD_i8_i8_2879_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2882_inst
    process(mul_val7_3_2684, mul_val8_3_2690) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_3_2684, mul_val8_3_2690, tmp_var);
      ADD_i8_i8_2882_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2883_inst
    process(ADD_i8_i8_2879_wire, ADD_i8_i8_2882_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2879_wire, ADD_i8_i8_2882_wire, tmp_var);
      ADD_i8_i8_2883_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2884_inst
    process(ADD_i8_i8_2876_wire, ADD_i8_i8_2883_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2876_wire, ADD_i8_i8_2883_wire, tmp_var);
      t_acc_val3_2885 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2889_inst
    process(mul_val1_4_2696, mul_val2_4_2702) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_4_2696, mul_val2_4_2702, tmp_var);
      ADD_i8_i8_2889_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2892_inst
    process(mul_val3_4_2708, mul_val4_4_2714) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_4_2708, mul_val4_4_2714, tmp_var);
      ADD_i8_i8_2892_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2893_inst
    process(ADD_i8_i8_2889_wire, ADD_i8_i8_2892_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2889_wire, ADD_i8_i8_2892_wire, tmp_var);
      ADD_i8_i8_2893_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2896_inst
    process(mul_val5_4_2720, mul_val6_4_2726) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_4_2720, mul_val6_4_2726, tmp_var);
      ADD_i8_i8_2896_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2899_inst
    process(mul_val7_4_2732, mul_val8_4_2738) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_4_2732, mul_val8_4_2738, tmp_var);
      ADD_i8_i8_2899_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2900_inst
    process(ADD_i8_i8_2896_wire, ADD_i8_i8_2899_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2896_wire, ADD_i8_i8_2899_wire, tmp_var);
      ADD_i8_i8_2900_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2901_inst
    process(ADD_i8_i8_2893_wire, ADD_i8_i8_2900_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2893_wire, ADD_i8_i8_2900_wire, tmp_var);
      t_acc_val4_2902 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2906_inst
    process(mul_val1_5_2744, mul_val2_5_2750) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_5_2744, mul_val2_5_2750, tmp_var);
      ADD_i8_i8_2906_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2909_inst
    process(mul_val3_5_2756, mul_val4_5_2762) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_5_2756, mul_val4_5_2762, tmp_var);
      ADD_i8_i8_2909_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2910_inst
    process(ADD_i8_i8_2906_wire, ADD_i8_i8_2909_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2906_wire, ADD_i8_i8_2909_wire, tmp_var);
      ADD_i8_i8_2910_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2913_inst
    process(mul_val5_5_2768, mul_val6_5_2774) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_5_2768, mul_val6_5_2774, tmp_var);
      ADD_i8_i8_2913_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2916_inst
    process(mul_val7_5_2780, mul_val8_5_2786) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_5_2780, mul_val8_5_2786, tmp_var);
      ADD_i8_i8_2916_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2917_inst
    process(ADD_i8_i8_2913_wire, ADD_i8_i8_2916_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2913_wire, ADD_i8_i8_2916_wire, tmp_var);
      ADD_i8_i8_2917_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2918_inst
    process(ADD_i8_i8_2910_wire, ADD_i8_i8_2917_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2910_wire, ADD_i8_i8_2917_wire, tmp_var);
      t_acc_val5_2919 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2923_inst
    process(mul_val1_6_2792, mul_val2_6_2798) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val1_6_2792, mul_val2_6_2798, tmp_var);
      ADD_i8_i8_2923_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2926_inst
    process(mul_val3_6_2804, mul_val4_6_2810) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val3_6_2804, mul_val4_6_2810, tmp_var);
      ADD_i8_i8_2926_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2927_inst
    process(ADD_i8_i8_2923_wire, ADD_i8_i8_2926_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2923_wire, ADD_i8_i8_2926_wire, tmp_var);
      ADD_i8_i8_2927_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2930_inst
    process(mul_val5_6_2816, mul_val6_6_2822) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val5_6_2816, mul_val6_6_2822, tmp_var);
      ADD_i8_i8_2930_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2933_inst
    process(mul_val7_6_2828, mul_val8_6_2834) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_val7_6_2828, mul_val8_6_2834, tmp_var);
      ADD_i8_i8_2933_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2934_inst
    process(ADD_i8_i8_2930_wire, ADD_i8_i8_2933_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2930_wire, ADD_i8_i8_2933_wire, tmp_var);
      ADD_i8_i8_2934_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2935_inst
    process(ADD_i8_i8_2927_wire, ADD_i8_i8_2934_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2927_wire, ADD_i8_i8_2934_wire, tmp_var);
      t_acc_val6_2936 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2943_inst
    process(acc1_2884_delayed_2_0_2939, t_acc_val1_2851) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc1_2884_delayed_2_0_2939, t_acc_val1_2851, tmp_var);
      ADD_i8_i8_2943_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2946_inst
    process(t_acc_val2_2868, t_acc_val3_2885) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(t_acc_val2_2868, t_acc_val3_2885, tmp_var);
      ADD_i8_i8_2946_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2947_inst
    process(ADD_i8_i8_2943_wire, ADD_i8_i8_2946_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2943_wire, ADD_i8_i8_2946_wire, tmp_var);
      acc_val1_2948 <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2955_inst
    process(acc2_2893_delayed_2_0_2951, t_acc_val4_2902) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(acc2_2893_delayed_2_0_2951, t_acc_val4_2902, tmp_var);
      ADD_i8_i8_2955_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2958_inst
    process(t_acc_val5_2919, t_acc_val6_2936) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(t_acc_val5_2919, t_acc_val6_2936, tmp_var);
      ADD_i8_i8_2958_wire <= tmp_var; --
    end process;
    -- binary operator ADD_i8_i8_2959_inst
    process(ADD_i8_i8_2955_wire, ADD_i8_i8_2958_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ADD_i8_i8_2955_wire, ADD_i8_i8_2958_wire, tmp_var);
      acc_val2_2960 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3030_inst
    process(chl_1919) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_1919, konst_3029_wire_constant, tmp_var);
      ADD_u16_u16_3030_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3050_inst
    process(col_1908) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_1908, konst_3049_wire_constant, tmp_var);
      ADD_u16_u16_3050_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3059_inst
    process(row_1903) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_1903, konst_3058_wire_constant, tmp_var);
      ADD_u16_u16_3059_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u2_u2_3039_inst
    process(num_1913) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_1913, konst_3038_wire_constant, tmp_var);
      ADD_u2_u2_3039_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2009_inst
    process(ULT_u16_u1_2005_wire, UGT_u2_u1_2008_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ULT_u16_u1_2005_wire, UGT_u2_u1_2008_wire, tmp_var);
      write_input_2010 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2302_inst
    process(EQ_u16_u1_2298_wire, EQ_u16_u1_2301_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u16_u1_2298_wire, EQ_u16_u1_2301_wire, tmp_var);
      read_k_2303 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2971_inst
    process(EQ_u2_u1_2969_wire, chl_done_2965) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_2969_wire, chl_done_2965, tmp_var);
      num_done_2972 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2981_inst
    process(col_done_2977, num_done_2972) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(col_done_2977, num_done_2972, tmp_var);
      row_done_2982 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2996_inst
    process(out_done_flag_2992, col_done_2977) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2992, col_done_2977, tmp_var);
      AND_u1_u1_2996_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3002_inst
    process(out_done_flag_2992, row_done_2982) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(out_done_flag_2992, row_done_2982, tmp_var);
      all_done_flag_3003 <= tmp_var; --
    end process;
    -- shared split operator group (58) : CONCAT_u8_u16_3090_inst 
    ApConcat_group_58: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3087_wire & type_cast_3089_wire;
      CONCAT_u8_u16_3090_wire <= data_out(15 downto 0);
      guard_vector(0)  <= num_done_3003_delayed_2_0_3083(0);
      reqL_unguarded(0) <= CONCAT_u8_u16_3090_inst_req_0;
      CONCAT_u8_u16_3090_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u8_u16_3090_inst_req_1;
      CONCAT_u8_u16_3090_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_58_gI: SplitGuardInterface generic map(name => "ApConcat_group_58_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_58",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- binary operator EQ_u16_u1_1928_inst
    process(col_1908) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1908, konst_1927_wire_constant, tmp_var);
      EQ_u16_u1_1928_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2298_inst
    process(col_1908) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1908, konst_2297_wire_constant, tmp_var);
      EQ_u16_u1_2298_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2301_inst
    process(row_1903) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(row_1903, konst_2300_wire_constant, tmp_var);
      EQ_u16_u1_2301_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2964_inst
    process(chl_1919, num_chl_1889) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(chl_1919, num_chl_1889, tmp_var);
      chl_done_2965 <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_2976_inst
    process(col_1908, num_col_1884) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_1908, num_col_1884, tmp_var);
      col_done_2977 <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1931_inst
    process(num_1913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_1913, konst_1930_wire_constant, tmp_var);
      EQ_u2_u1_1931_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_2969_inst
    process(num_1913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(num_1913, konst_2968_wire_constant, tmp_var);
      EQ_u2_u1_2969_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2550_inst
    process(kval1_1_2454, ival1_1_2170) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_1_2454, ival1_1_2170, tmp_var);
      MUL_i8_i8_2550_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2556_inst
    process(kval2_1_2458, ival2_1_2174) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_1_2458, ival2_1_2174, tmp_var);
      MUL_i8_i8_2556_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2562_inst
    process(kval3_1_2462, ival3_1_2178) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_1_2462, ival3_1_2178, tmp_var);
      MUL_i8_i8_2562_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2568_inst
    process(kval4_1_2466, ival4_1_2182) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_1_2466, ival4_1_2182, tmp_var);
      MUL_i8_i8_2568_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2574_inst
    process(kval5_1_2470, ival5_1_2186) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_1_2470, ival5_1_2186, tmp_var);
      MUL_i8_i8_2574_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2580_inst
    process(kval6_1_2474, ival6_1_2190) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_1_2474, ival6_1_2190, tmp_var);
      MUL_i8_i8_2580_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2586_inst
    process(kval7_1_2478, ival7_1_2194) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_1_2478, ival7_1_2194, tmp_var);
      MUL_i8_i8_2586_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2592_inst
    process(kval8_1_2482, ival8_1_2198) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_1_2482, ival8_1_2198, tmp_var);
      MUL_i8_i8_2592_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2598_inst
    process(kval1_2_2486, ival1_2_2202) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2_2486, ival1_2_2202, tmp_var);
      MUL_i8_i8_2598_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2604_inst
    process(kval2_2_2490, ival2_2_2206) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2_2490, ival2_2_2206, tmp_var);
      MUL_i8_i8_2604_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2610_inst
    process(kval3_2_2494, ival3_2_2210) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2_2494, ival3_2_2210, tmp_var);
      MUL_i8_i8_2610_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2616_inst
    process(kval4_2_2498, ival4_2_2214) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_2_2498, ival4_2_2214, tmp_var);
      MUL_i8_i8_2616_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2622_inst
    process(kval5_2_2502, ival5_2_2218) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_2_2502, ival5_2_2218, tmp_var);
      MUL_i8_i8_2622_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2628_inst
    process(kval6_2_2506, ival6_2_2222) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_2_2506, ival6_2_2222, tmp_var);
      MUL_i8_i8_2628_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2634_inst
    process(kval7_2_2510, ival7_2_2226) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_2_2510, ival7_2_2226, tmp_var);
      MUL_i8_i8_2634_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2640_inst
    process(kval8_2_2514, ival8_2_2230) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_2_2514, ival8_2_2230, tmp_var);
      MUL_i8_i8_2640_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2646_inst
    process(kval1_3_2518, ival1_3_2234) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_3_2518, ival1_3_2234, tmp_var);
      MUL_i8_i8_2646_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2652_inst
    process(kval2_3_2522, ival2_3_2238) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_3_2522, ival2_3_2238, tmp_var);
      MUL_i8_i8_2652_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2658_inst
    process(kval3_3_2526, ival3_3_2242) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_3_2526, ival3_3_2242, tmp_var);
      MUL_i8_i8_2658_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2664_inst
    process(kval4_3_2530, ival4_3_2246) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_3_2530, ival4_3_2246, tmp_var);
      MUL_i8_i8_2664_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2670_inst
    process(kval5_3_2534, ival5_3_2250) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_3_2534, ival5_3_2250, tmp_var);
      MUL_i8_i8_2670_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2676_inst
    process(kval6_3_2538, ival6_3_2254) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_3_2538, ival6_3_2254, tmp_var);
      MUL_i8_i8_2676_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2682_inst
    process(kval7_3_2542, ival7_3_2258) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_3_2542, ival7_3_2258, tmp_var);
      MUL_i8_i8_2682_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2688_inst
    process(kval8_3_2546, ival8_3_2262) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_3_2546, ival8_3_2262, tmp_var);
      MUL_i8_i8_2688_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2694_inst
    process(kval1_1_2454, ival1_2_2202) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_1_2454, ival1_2_2202, tmp_var);
      MUL_i8_i8_2694_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2700_inst
    process(kval2_1_2458, ival2_2_2206) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_1_2458, ival2_2_2206, tmp_var);
      MUL_i8_i8_2700_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2706_inst
    process(kval3_1_2462, ival3_2_2210) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_1_2462, ival3_2_2210, tmp_var);
      MUL_i8_i8_2706_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2712_inst
    process(kval4_1_2466, ival4_2_2214) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_1_2466, ival4_2_2214, tmp_var);
      MUL_i8_i8_2712_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2718_inst
    process(kval5_1_2470, ival5_2_2218) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_1_2470, ival5_2_2218, tmp_var);
      MUL_i8_i8_2718_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2724_inst
    process(kval6_1_2474, ival6_2_2222) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_1_2474, ival6_2_2222, tmp_var);
      MUL_i8_i8_2724_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2730_inst
    process(kval7_1_2478, ival7_2_2226) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_1_2478, ival7_2_2226, tmp_var);
      MUL_i8_i8_2730_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2736_inst
    process(kval8_1_2482, ival8_2_2230) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_1_2482, ival8_2_2230, tmp_var);
      MUL_i8_i8_2736_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2742_inst
    process(kval1_2_2486, ival1_3_2234) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_2_2486, ival1_3_2234, tmp_var);
      MUL_i8_i8_2742_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2748_inst
    process(kval2_2_2490, ival2_3_2238) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_2_2490, ival2_3_2238, tmp_var);
      MUL_i8_i8_2748_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2754_inst
    process(kval3_2_2494, ival3_3_2242) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_2_2494, ival3_3_2242, tmp_var);
      MUL_i8_i8_2754_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2760_inst
    process(kval4_2_2498, ival4_3_2246) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_2_2498, ival4_3_2246, tmp_var);
      MUL_i8_i8_2760_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2766_inst
    process(kval5_2_2502, ival5_3_2250) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_2_2502, ival5_3_2250, tmp_var);
      MUL_i8_i8_2766_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2772_inst
    process(kval6_2_2506, ival6_3_2254) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_2_2506, ival6_3_2254, tmp_var);
      MUL_i8_i8_2772_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2778_inst
    process(kval7_2_2510, ival7_3_2258) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_2_2510, ival7_3_2258, tmp_var);
      MUL_i8_i8_2778_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2784_inst
    process(kval8_2_2514, ival8_3_2262) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_2_2514, ival8_3_2262, tmp_var);
      MUL_i8_i8_2784_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2790_inst
    process(kval1_3_2518, ival1_4_2266) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval1_3_2518, ival1_4_2266, tmp_var);
      MUL_i8_i8_2790_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2796_inst
    process(kval2_3_2522, ival2_4_2270) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval2_3_2522, ival2_4_2270, tmp_var);
      MUL_i8_i8_2796_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2802_inst
    process(kval3_3_2526, ival3_4_2274) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval3_3_2526, ival3_4_2274, tmp_var);
      MUL_i8_i8_2802_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2808_inst
    process(kval4_3_2530, ival4_4_2278) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval4_3_2530, ival4_4_2278, tmp_var);
      MUL_i8_i8_2808_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2814_inst
    process(kval5_3_2534, ival5_4_2282) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval5_3_2534, ival5_4_2282, tmp_var);
      MUL_i8_i8_2814_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2820_inst
    process(kval6_3_2538, ival6_4_2286) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval6_3_2538, ival6_4_2286, tmp_var);
      MUL_i8_i8_2820_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2826_inst
    process(kval7_3_2542, ival7_4_2290) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval7_3_2542, ival7_4_2290, tmp_var);
      MUL_i8_i8_2826_wire <= tmp_var; --
    end process;
    -- binary operator MUL_i8_i8_2832_inst
    process(kval8_3_2546, ival8_4_2294) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntMul_proc(kval8_3_2546, ival8_4_2294, tmp_var);
      MUL_i8_i8_2832_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2997_inst
    process(AND_u1_u1_2996_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", AND_u1_u1_2996_wire, tmp_var);
      store_kernel_2998 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3094_inst
    process(all_done_flag_3003) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", all_done_flag_3003, tmp_var);
      NOT_u1_u1_3094_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1932_inst
    process(EQ_u16_u1_1928_wire, EQ_u2_u1_1931_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u16_u1_1928_wire, EQ_u2_u1_1931_wire, tmp_var);
      read_ip_1933 <= tmp_var; --
    end process;
    -- shared split operator group (117) : SUB_u16_u16_1878_inst 
    ApIntSub_group_117: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_1876_wire;
      num_row_1879 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1878_inst_req_0;
      SUB_u16_u16_1878_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1878_inst_req_1;
      SUB_u16_u16_1878_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_117_gI: SplitGuardInterface generic map(name => "ApIntSub_group_117_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_117",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 117
    -- shared split operator group (118) : SUB_u16_u16_1883_inst 
    ApIntSub_group_118: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_num_out_pipe_1881_wire;
      num_col_1884 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1883_inst_req_0;
      SUB_u16_u16_1883_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1883_inst_req_1;
      SUB_u16_u16_1883_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_118_gI: SplitGuardInterface generic map(name => "ApIntSub_group_118_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_118",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 118
    -- shared split operator group (119) : SUB_u16_u16_1888_inst 
    ApIntSub_group_119: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= RPIPE_size_pipe_1886_wire;
      num_chl_1889 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_1888_inst_req_0;
      SUB_u16_u16_1888_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_1888_inst_req_1;
      SUB_u16_u16_1888_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_119_gI: SplitGuardInterface generic map(name => "ApIntSub_group_119_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_119",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 119
    -- shared split operator group (120) : SUB_u16_u16_2986_inst 
    ApIntSub_group_120: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= num_row_1879;
      SUB_u16_u16_2927_2927_delayed_1_0_2987 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_2986_inst_req_0;
      SUB_u16_u16_2986_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_2986_inst_req_1;
      SUB_u16_u16_2986_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_120_gI: SplitGuardInterface generic map(name => "ApIntSub_group_120_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_120",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 120
    -- binary operator UGE_u16_u1_2991_inst
    process(row_1903, SUB_u16_u16_2927_2927_delayed_1_0_2987) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_1903, SUB_u16_u16_2927_2927_delayed_1_0_2987, tmp_var);
      out_done_flag_2992 <= tmp_var; --
    end process;
    -- binary operator UGT_u2_u1_2008_inst
    process(num_1913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(num_1913, konst_2007_wire_constant, tmp_var);
      UGT_u2_u1_2008_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_2005_inst
    process(col_1908, num_col_1884) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(col_1908, num_col_1884, tmp_var);
      ULT_u16_u1_2005_wire <= tmp_var; --
    end process;
    xxconvolvexxconv_ip1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip1",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip1_pipe_read_req,
        read_ack => xxconvolvexxconv_ip1_pipe_read_ack,
        read_data => xxconvolvexxconv_ip1_pipe_read_data,
        write_req => xxconvolvexxconv_ip1_pipe_write_req,
        write_ack => xxconvolvexxconv_ip1_pipe_write_ack,
        write_data => xxconvolvexxconv_ip1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip2",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip2_pipe_read_req,
        read_ack => xxconvolvexxconv_ip2_pipe_read_ack,
        read_data => xxconvolvexxconv_ip2_pipe_read_data,
        write_req => xxconvolvexxconv_ip2_pipe_write_req,
        write_ack => xxconvolvexxconv_ip2_pipe_write_ack,
        write_data => xxconvolvexxconv_ip2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip3",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip3_pipe_read_req,
        read_ack => xxconvolvexxconv_ip3_pipe_read_ack,
        read_data => xxconvolvexxconv_ip3_pipe_read_data,
        write_req => xxconvolvexxconv_ip3_pipe_write_req,
        write_ack => xxconvolvexxconv_ip3_pipe_write_ack,
        write_data => xxconvolvexxconv_ip3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_ip4_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_ip4",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_ip4_pipe_read_req,
        read_ack => xxconvolvexxconv_ip4_pipe_read_ack,
        read_data => xxconvolvexxconv_ip4_pipe_read_data,
        write_req => xxconvolvexxconv_ip4_pipe_write_req,
        write_ack => xxconvolvexxconv_ip4_pipe_write_ack,
        write_data => xxconvolvexxconv_ip4_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k1_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k1",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k1_pipe_read_req,
        read_ack => xxconvolvexxconv_k1_pipe_read_ack,
        read_data => xxconvolvexxconv_k1_pipe_read_data,
        write_req => xxconvolvexxconv_k1_pipe_write_req,
        write_ack => xxconvolvexxconv_k1_pipe_write_ack,
        write_data => xxconvolvexxconv_k1_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k2_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k2",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k2_pipe_read_req,
        read_ack => xxconvolvexxconv_k2_pipe_read_ack,
        read_data => xxconvolvexxconv_k2_pipe_read_data,
        write_req => xxconvolvexxconv_k2_pipe_write_req,
        write_ack => xxconvolvexxconv_k2_pipe_write_ack,
        write_data => xxconvolvexxconv_k2_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxconvolvexxconv_k3_Pipe: PipeBase -- 
      generic map( -- 
        name => "pipe xxconvolvexxconv_k3",
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        lifo_mode => false,
        full_rate => false,
        shift_register_mode => false,
        bypass => false,
        depth => 512 --
      )
      port map( -- 
        read_req => xxconvolvexxconv_k3_pipe_read_req,
        read_ack => xxconvolvexxconv_k3_pipe_read_ack,
        read_data => xxconvolvexxconv_k3_pipe_read_data,
        write_req => xxconvolvexxconv_k3_pipe_write_req,
        write_ack => xxconvolvexxconv_k3_pipe_write_ack,
        write_data => xxconvolvexxconv_k3_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : RPIPE_input_pipe1_1936_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe1_1936_inst_req_0;
      RPIPE_input_pipe1_1936_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe1_1936_inst_req_1;
      RPIPE_input_pipe1_1936_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1933(0);
      temp2_1_1937 <= data_out(63 downto 0);
      input_pipe1_read_0_gI: SplitGuardInterface generic map(name => "input_pipe1_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe1_read_0: InputPortRevised -- 
        generic map ( name => "input_pipe1_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe1_pipe_read_req(0),
          oack => input_pipe1_pipe_read_ack(0),
          odata => input_pipe1_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_input_pipe2_1940_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe2_1940_inst_req_0;
      RPIPE_input_pipe2_1940_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe2_1940_inst_req_1;
      RPIPE_input_pipe2_1940_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1933(0);
      temp2_2_1941 <= data_out(63 downto 0);
      input_pipe2_read_1_gI: SplitGuardInterface generic map(name => "input_pipe2_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe2_read_1: InputPortRevised -- 
        generic map ( name => "input_pipe2_read_1", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe2_pipe_read_req(0),
          oack => input_pipe2_pipe_read_ack(0),
          odata => input_pipe2_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_input_pipe3_1944_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe3_1944_inst_req_0;
      RPIPE_input_pipe3_1944_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe3_1944_inst_req_1;
      RPIPE_input_pipe3_1944_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1933(0);
      temp2_3_1945 <= data_out(63 downto 0);
      input_pipe3_read_2_gI: SplitGuardInterface generic map(name => "input_pipe3_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe3_read_2: InputPortRevised -- 
        generic map ( name => "input_pipe3_read_2", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe3_pipe_read_req(0),
          oack => input_pipe3_pipe_read_ack(0),
          odata => input_pipe3_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_input_pipe4_1948_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_pipe4_1948_inst_req_0;
      RPIPE_input_pipe4_1948_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_pipe4_1948_inst_req_1;
      RPIPE_input_pipe4_1948_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_ip_1933(0);
      temp2_4_1949 <= data_out(63 downto 0);
      input_pipe4_read_3_gI: SplitGuardInterface generic map(name => "input_pipe4_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_pipe4_read_3: InputPortRevised -- 
        generic map ( name => "input_pipe4_read_3", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_pipe4_pipe_read_req(0),
          oack => input_pipe4_pipe_read_ack(0),
          odata => input_pipe4_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : RPIPE_kernel_pipe1_2306_inst 
    InportGroup_4: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe1_2306_inst_req_0;
      RPIPE_kernel_pipe1_2306_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe1_2306_inst_req_1;
      RPIPE_kernel_pipe1_2306_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2303(0);
      tempk1_1_2307 <= data_out(63 downto 0);
      kernel_pipe1_read_4_gI: SplitGuardInterface generic map(name => "kernel_pipe1_read_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_read_4: InputPortRevised -- 
        generic map ( name => "kernel_pipe1_read_4", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe1_pipe_read_req(0),
          oack => kernel_pipe1_pipe_read_ack(0),
          odata => kernel_pipe1_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : RPIPE_kernel_pipe2_2310_inst 
    InportGroup_5: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe2_2310_inst_req_0;
      RPIPE_kernel_pipe2_2310_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe2_2310_inst_req_1;
      RPIPE_kernel_pipe2_2310_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2303(0);
      tempk1_2_2311 <= data_out(63 downto 0);
      kernel_pipe2_read_5_gI: SplitGuardInterface generic map(name => "kernel_pipe2_read_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_read_5: InputPortRevised -- 
        generic map ( name => "kernel_pipe2_read_5", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe2_pipe_read_req(0),
          oack => kernel_pipe2_pipe_read_ack(0),
          odata => kernel_pipe2_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : RPIPE_kernel_pipe3_2314_inst 
    InportGroup_6: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_kernel_pipe3_2314_inst_req_0;
      RPIPE_kernel_pipe3_2314_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_kernel_pipe3_2314_inst_req_1;
      RPIPE_kernel_pipe3_2314_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= read_k_2303(0);
      tempk1_3_2315 <= data_out(63 downto 0);
      kernel_pipe3_read_6_gI: SplitGuardInterface generic map(name => "kernel_pipe3_read_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_read_6: InputPortRevised -- 
        generic map ( name => "kernel_pipe3_read_6", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => kernel_pipe3_pipe_read_req(0),
          oack => kernel_pipe3_pipe_read_ack(0),
          odata => kernel_pipe3_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : RPIPE_num_out_pipe_1876_inst RPIPE_num_out_pipe_1881_inst 
    InportGroup_7: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 1 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= RPIPE_num_out_pipe_1876_inst_req_0;
      reqL_unguarded(0) <= RPIPE_num_out_pipe_1881_inst_req_0;
      RPIPE_num_out_pipe_1876_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_num_out_pipe_1881_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= RPIPE_num_out_pipe_1876_inst_req_1;
      reqR_unguarded(0) <= RPIPE_num_out_pipe_1881_inst_req_1;
      RPIPE_num_out_pipe_1876_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_num_out_pipe_1881_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      RPIPE_num_out_pipe_1876_wire <= data_out(31 downto 16);
      RPIPE_num_out_pipe_1881_wire <= data_out(15 downto 0);
      num_out_pipe_read_7_gI: SplitGuardInterface generic map(name => "num_out_pipe_read_7_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      num_out_pipe_read_7: InputPortRevised -- 
        generic map ( name => "num_out_pipe_read_7", data_width => 16,  num_reqs => 2,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => num_out_pipe_pipe_read_req(0),
          oack => num_out_pipe_pipe_read_ack(0),
          odata => num_out_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : RPIPE_size_pipe_1886_inst 
    InportGroup_8: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_size_pipe_1886_inst_req_0;
      RPIPE_size_pipe_1886_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_size_pipe_1886_inst_req_1;
      RPIPE_size_pipe_1886_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_size_pipe_1886_wire <= data_out(15 downto 0);
      size_pipe_read_8_gI: SplitGuardInterface generic map(name => "size_pipe_read_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      size_pipe_read_8: InputPortRevised -- 
        generic map ( name => "size_pipe_read_8", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => size_pipe_pipe_read_req(0),
          oack => size_pipe_pipe_read_ack(0),
          odata => size_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : RPIPE_xxconvolvexxconv_ip1_1952_inst 
    InportGroup_9: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_1952_inst_req_0;
      RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip1_1952_inst_req_1;
      RPIPE_xxconvolvexxconv_ip1_1952_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1933(0);
      temp1_1_1953 <= data_out(63 downto 0);
      xxconvolvexxconv_ip1_read_9_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_read_9_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_read_9: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1_read_9", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip1_pipe_read_req(0),
          oack => xxconvolvexxconv_ip1_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : RPIPE_xxconvolvexxconv_ip2_1956_inst 
    InportGroup_10: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_1956_inst_req_0;
      RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip2_1956_inst_req_1;
      RPIPE_xxconvolvexxconv_ip2_1956_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1933(0);
      temp1_2_1957 <= data_out(63 downto 0);
      xxconvolvexxconv_ip2_read_10_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_read_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_read_10: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2_read_10", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip2_pipe_read_req(0),
          oack => xxconvolvexxconv_ip2_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : RPIPE_xxconvolvexxconv_ip3_1960_inst 
    InportGroup_11: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_1960_inst_req_0;
      RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip3_1960_inst_req_1;
      RPIPE_xxconvolvexxconv_ip3_1960_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1933(0);
      temp1_3_1961 <= data_out(63 downto 0);
      xxconvolvexxconv_ip3_read_11_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_read_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_read_11: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3_read_11", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip3_pipe_read_req(0),
          oack => xxconvolvexxconv_ip3_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : RPIPE_xxconvolvexxconv_ip4_1964_inst 
    InportGroup_12: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_1964_inst_req_0;
      RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_ip4_1964_inst_req_1;
      RPIPE_xxconvolvexxconv_ip4_1964_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_ip_1933(0);
      temp1_4_1965 <= data_out(63 downto 0);
      xxconvolvexxconv_ip4_read_12_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_read_12_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_read_12: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4_read_12", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_ip4_pipe_read_req(0),
          oack => xxconvolvexxconv_ip4_pipe_read_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- shared inport operator group (13) : RPIPE_xxconvolvexxconv_k1_2318_inst 
    InportGroup_13: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2318_inst_req_0;
      RPIPE_xxconvolvexxconv_k1_2318_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k1_2318_inst_req_1;
      RPIPE_xxconvolvexxconv_k1_2318_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2303(0);
      tempk2_1_2319 <= data_out(63 downto 0);
      xxconvolvexxconv_k1_read_13_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_read_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_read_13: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1_read_13", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k1_pipe_read_req(0),
          oack => xxconvolvexxconv_k1_pipe_read_ack(0),
          odata => xxconvolvexxconv_k1_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 13
    -- shared inport operator group (14) : RPIPE_xxconvolvexxconv_k2_2322_inst 
    InportGroup_14: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2322_inst_req_0;
      RPIPE_xxconvolvexxconv_k2_2322_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k2_2322_inst_req_1;
      RPIPE_xxconvolvexxconv_k2_2322_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2303(0);
      tempk2_2_2323 <= data_out(63 downto 0);
      xxconvolvexxconv_k2_read_14_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_read_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_read_14: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2_read_14", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k2_pipe_read_req(0),
          oack => xxconvolvexxconv_k2_pipe_read_ack(0),
          odata => xxconvolvexxconv_k2_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 14
    -- shared inport operator group (15) : RPIPE_xxconvolvexxconv_k3_2326_inst 
    InportGroup_15: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2326_inst_req_0;
      RPIPE_xxconvolvexxconv_k3_2326_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_xxconvolvexxconv_k3_2326_inst_req_1;
      RPIPE_xxconvolvexxconv_k3_2326_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not read_k_2303(0);
      tempk2_3_2327 <= data_out(63 downto 0);
      xxconvolvexxconv_k3_read_15_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_read_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_read_15: InputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3_read_15", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => xxconvolvexxconv_k3_pipe_read_req(0),
          oack => xxconvolvexxconv_k3_pipe_read_ack(0),
          odata => xxconvolvexxconv_k3_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 15
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3095_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3095_inst_req_0;
      WPIPE_input_done_pipe_3095_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3095_inst_req_1;
      WPIPE_input_done_pipe_3095_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3096_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_output_pipe_3085_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_output_pipe_3085_inst_req_0;
      WPIPE_output_pipe_3085_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_output_pipe_3085_inst_req_1;
      WPIPE_output_pipe_3085_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= num_done_3003_delayed_2_0_3083(0);
      data_in <= CONCAT_u8_u16_3090_wire;
      output_pipe_write_1_gI: SplitGuardInterface generic map(name => "output_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      output_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "output_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => output_pipe_pipe_write_req(0),
          oack => output_pipe_pipe_write_ack(0),
          odata => output_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_xxconvolvexxconv_ip1_2015_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2015_inst_req_0;
      WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip1_2015_inst_req_1;
      WPIPE_xxconvolvexxconv_ip1_2015_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1978_delayed_1_0_2013(0);
      data_in <= iread1_1974;
      xxconvolvexxconv_ip1_write_2_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip1_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip1_write_2: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip1", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip1_pipe_write_req(0),
          oack => xxconvolvexxconv_ip1_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip1_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_xxconvolvexxconv_ip2_2022_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2022_inst_req_0;
      WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip2_2022_inst_req_1;
      WPIPE_xxconvolvexxconv_ip2_2022_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1982_delayed_1_0_2020(0);
      data_in <= iread2_1983;
      xxconvolvexxconv_ip2_write_3_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip2_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip2_write_3: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip2", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip2_pipe_write_req(0),
          oack => xxconvolvexxconv_ip2_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip2_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_xxconvolvexxconv_ip3_2029_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2029_inst_req_0;
      WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip3_2029_inst_req_1;
      WPIPE_xxconvolvexxconv_ip3_2029_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1986_delayed_1_0_2027(0);
      data_in <= iread3_1992;
      xxconvolvexxconv_ip3_write_4_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip3_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip3_write_4: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip3", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip3_pipe_write_req(0),
          oack => xxconvolvexxconv_ip3_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip3_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared outport operator group (5) : WPIPE_xxconvolvexxconv_ip4_2036_inst 
    OutportGroup_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2036_inst_req_0;
      WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_ip4_2036_inst_req_1;
      WPIPE_xxconvolvexxconv_ip4_2036_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_input_1990_delayed_1_0_2034(0);
      data_in <= iread4_2001;
      xxconvolvexxconv_ip4_write_5_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_ip4_write_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_ip4_write_5: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_ip4", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_ip4_pipe_write_req(0),
          oack => xxconvolvexxconv_ip4_pipe_write_ack(0),
          odata => xxconvolvexxconv_ip4_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- shared outport operator group (6) : WPIPE_xxconvolvexxconv_k1_3008_inst 
    OutportGroup_6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_3008_inst_req_0;
      WPIPE_xxconvolvexxconv_k1_3008_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k1_3008_inst_req_1;
      WPIPE_xxconvolvexxconv_k1_3008_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2941_delayed_1_0_3006(0);
      data_in <= kread1_2336;
      xxconvolvexxconv_k1_write_6_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k1_write_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k1_write_6: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k1", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k1_pipe_write_req(0),
          oack => xxconvolvexxconv_k1_pipe_write_ack(0),
          odata => xxconvolvexxconv_k1_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- shared outport operator group (7) : WPIPE_xxconvolvexxconv_k2_3015_inst 
    OutportGroup_7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_3015_inst_req_0;
      WPIPE_xxconvolvexxconv_k2_3015_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k2_3015_inst_req_1;
      WPIPE_xxconvolvexxconv_k2_3015_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2945_delayed_1_0_3013(0);
      data_in <= kread2_2345;
      xxconvolvexxconv_k2_write_7_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k2_write_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k2_write_7: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k2", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k2_pipe_write_req(0),
          oack => xxconvolvexxconv_k2_pipe_write_ack(0),
          odata => xxconvolvexxconv_k2_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- shared outport operator group (8) : WPIPE_xxconvolvexxconv_k3_3022_inst 
    OutportGroup_8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_3022_inst_req_0;
      WPIPE_xxconvolvexxconv_k3_3022_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_xxconvolvexxconv_k3_3022_inst_req_1;
      WPIPE_xxconvolvexxconv_k3_3022_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= store_kernel_2949_delayed_1_0_3020(0);
      data_in <= kread3_2354;
      xxconvolvexxconv_k3_write_8_gI: SplitGuardInterface generic map(name => "xxconvolvexxconv_k3_write_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      xxconvolvexxconv_k3_write_8: OutputPortRevised -- 
        generic map ( name => "xxconvolvexxconv_k3", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => xxconvolvexxconv_k3_pipe_write_req(0),
          oack => xxconvolvexxconv_k3_pipe_write_ack(0),
          odata => xxconvolvexxconv_k3_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- 
  end Block; -- data_path
  -- 
end convolve_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity loadKernelChannel is -- 
  generic (tag_length : integer); 
  port ( -- 
    start_add : in  std_logic_vector(31 downto 0);
    num_chl : in  std_logic_vector(15 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
    input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
    kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
    kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
    kernel_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
    size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadKernelChannel;
architecture loadKernelChannel_arch of loadKernelChannel is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 48)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal start_add_buffer :  std_logic_vector(31 downto 0);
  signal start_add_update_enable: Boolean;
  signal num_chl_buffer :  std_logic_vector(15 downto 0);
  signal num_chl_update_enable: Boolean;
  -- output port buffer signals
  signal loadKernelChannel_CP_1349_start: Boolean;
  signal loadKernelChannel_CP_1349_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal addr_of_469_final_reg_req_1 : boolean;
  signal start_add_456_buf_req_0 : boolean;
  signal addr_of_469_final_reg_ack_1 : boolean;
  signal nmycount_462_455_buf_ack_0 : boolean;
  signal nmycount_462_455_buf_req_0 : boolean;
  signal addr_of_469_final_reg_ack_0 : boolean;
  signal array_obj_ref_468_index_offset_ack_1 : boolean;
  signal array_obj_ref_468_index_offset_req_1 : boolean;
  signal addr_of_469_final_reg_req_0 : boolean;
  signal array_obj_ref_468_index_offset_req_0 : boolean;
  signal start_add_456_buf_req_1 : boolean;
  signal RPIPE_input_done_pipe_448_inst_ack_1 : boolean;
  signal start_add_456_buf_ack_0 : boolean;
  signal W_send_to_1_481_delayed_13_0_493_inst_req_0 : boolean;
  signal ptr_deref_473_load_0_req_0 : boolean;
  signal start_add_456_buf_ack_1 : boolean;
  signal nmycount_462_455_buf_req_1 : boolean;
  signal nmycount_462_455_buf_ack_1 : boolean;
  signal do_while_stmt_451_branch_req_0 : boolean;
  signal phi_stmt_453_req_0 : boolean;
  signal phi_stmt_453_req_1 : boolean;
  signal ptr_deref_473_load_0_ack_0 : boolean;
  signal W_send_to_1_481_delayed_13_0_493_inst_ack_0 : boolean;
  signal W_send_to_1_481_delayed_13_0_493_inst_req_1 : boolean;
  signal phi_stmt_453_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_ack_1 : boolean;
  signal ptr_deref_473_load_0_req_1 : boolean;
  signal W_send_to_1_481_delayed_13_0_493_inst_ack_1 : boolean;
  signal ptr_deref_473_load_0_ack_1 : boolean;
  signal RPIPE_input_done_pipe_448_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_ack_0 : boolean;
  signal W_send_to_2_485_delayed_13_0_500_inst_req_1 : boolean;
  signal array_obj_ref_468_index_offset_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_504_inst_ack_1 : boolean;
  signal RPIPE_input_done_pipe_448_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe1_497_inst_req_1 : boolean;
  signal RPIPE_input_done_pipe_448_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe2_504_inst_req_0 : boolean;
  signal W_send_to_2_485_delayed_13_0_500_inst_ack_1 : boolean;
  signal W_send_to_2_485_delayed_13_0_500_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_504_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe2_504_inst_req_1 : boolean;
  signal W_send_to_3_489_delayed_13_0_507_inst_req_1 : boolean;
  signal W_send_to_3_489_delayed_13_0_507_inst_ack_1 : boolean;
  signal W_send_to_2_485_delayed_13_0_500_inst_req_0 : boolean;
  signal W_send_to_3_489_delayed_13_0_507_inst_req_0 : boolean;
  signal W_send_to_3_489_delayed_13_0_507_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_511_inst_req_0 : boolean;
  signal WPIPE_kernel_pipe3_511_inst_ack_0 : boolean;
  signal WPIPE_kernel_pipe3_511_inst_req_1 : boolean;
  signal WPIPE_kernel_pipe3_511_inst_ack_1 : boolean;
  signal do_while_stmt_451_branch_ack_0 : boolean;
  signal do_while_stmt_451_branch_ack_1 : boolean;
  signal WPIPE_size_pipe_521_inst_req_0 : boolean;
  signal WPIPE_size_pipe_521_inst_ack_0 : boolean;
  signal WPIPE_size_pipe_521_inst_req_1 : boolean;
  signal WPIPE_size_pipe_521_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadKernelChannel_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 48) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= start_add;
  start_add_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(47 downto 32) <= num_chl;
  num_chl_buffer <= in_buffer_data_out(47 downto 32);
  in_buffer_data_in(tag_length + 47 downto 48) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 47 downto 48);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadKernelChannel_CP_1349_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadKernelChannel_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1349_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1349_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadKernelChannel_CP_1349_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadKernelChannel_CP_1349: Block -- control-path 
    signal loadKernelChannel_CP_1349_elements: BooleanArray(69 downto 0);
    -- 
  begin -- 
    loadKernelChannel_CP_1349_elements(0) <= loadKernelChannel_CP_1349_start;
    loadKernelChannel_CP_1349_symbol <= loadKernelChannel_CP_1349_elements(69);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_420_to_assign_stmt_449/$entry
      -- CP-element group 0: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Sample/rr
      -- CP-element group 0: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_sample_start_
      -- 
    rr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(0), ack => RPIPE_input_done_pipe_448_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Update/cr
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Update/$entry
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Sample/ra
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_update_start_
      -- CP-element group 1: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_sample_completed_
      -- 
    ra_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_448_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(1)); -- 
    cr_1367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(1), ack => RPIPE_input_done_pipe_448_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 branch_block_stmt_450/$entry
      -- CP-element group 2: 	 branch_block_stmt_450/do_while_stmt_451__entry__
      -- CP-element group 2: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_450/branch_block_stmt_450__entry__
      -- CP-element group 2: 	 assign_stmt_420_to_assign_stmt_449/$exit
      -- CP-element group 2: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_Update/$exit
      -- CP-element group 2: 	 assign_stmt_420_to_assign_stmt_449/RPIPE_input_done_pipe_448_update_completed_
      -- 
    ca_1368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_input_done_pipe_448_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(2)); -- 
    -- CP-element group 3:  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	67 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	68 
    -- CP-element group 3:  members (7) 
      -- CP-element group 3: 	 branch_block_stmt_450/branch_block_stmt_450__exit__
      -- CP-element group 3: 	 branch_block_stmt_450/do_while_stmt_451__exit__
      -- CP-element group 3: 	 branch_block_stmt_450/$exit
      -- CP-element group 3: 	 assign_stmt_523/$entry
      -- CP-element group 3: 	 assign_stmt_523/WPIPE_size_pipe_521_sample_start_
      -- CP-element group 3: 	 assign_stmt_523/WPIPE_size_pipe_521_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_523/WPIPE_size_pipe_521_Sample/req
      -- 
    req_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(3), ack => WPIPE_size_pipe_521_inst_req_0); -- 
    loadKernelChannel_CP_1349_elements(3) <= loadKernelChannel_CP_1349_elements(67);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_450/do_while_stmt_451/$entry
      -- CP-element group 4: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451__entry__
      -- 
    loadKernelChannel_CP_1349_elements(4) <= loadKernelChannel_CP_1349_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	67 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451__exit__
      -- 
    -- Element group loadKernelChannel_CP_1349_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_450/do_while_stmt_451/loop_back
      -- 
    -- Element group loadKernelChannel_CP_1349_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	65 
    -- CP-element group 7: 	66 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_450/do_while_stmt_451/condition_done
      -- CP-element group 7: 	 branch_block_stmt_450/do_while_stmt_451/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_450/do_while_stmt_451/loop_taken/$entry
      -- 
    loadKernelChannel_CP_1349_elements(7) <= loadKernelChannel_CP_1349_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	64 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_450/do_while_stmt_451/loop_body_done
      -- 
    loadKernelChannel_CP_1349_elements(8) <= loadKernelChannel_CP_1349_elements(64);
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	18 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/back_edge_to_loop_body
      -- 
    loadKernelChannel_CP_1349_elements(9) <= loadKernelChannel_CP_1349_elements(6);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	20 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/first_time_through_loop_body
      -- 
    loadKernelChannel_CP_1349_elements(10) <= loadKernelChannel_CP_1349_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	32 
    -- CP-element group 11: 	33 
    -- CP-element group 11: 	63 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/loop_body_start
      -- 
    -- Element group loadKernelChannel_CP_1349_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	63 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/condition_evaluated
      -- 
    condition_evaluated_1390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(12), ack => do_while_stmt_451_branch_req_0); -- 
    loadKernelChannel_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(17) & loadKernelChannel_CP_1349_elements(63);
      gj_loadKernelChannel_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/aggregated_phi_sample_req
      -- 
    loadKernelChannel_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(14) & loadKernelChannel_CP_1349_elements(17);
      gj_loadKernelChannel_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	13 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_sample_start_
      -- 
    loadKernelChannel_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(11) & loadKernelChannel_CP_1349_elements(16);
      gj_loadKernelChannel_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	34 
    -- CP-element group 15: 	44 
    -- CP-element group 15: 	51 
    -- CP-element group 15: 	58 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_update_start_
      -- CP-element group 15: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_update_start__ps
      -- CP-element group 15: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/aggregated_phi_update_req
      -- 
    loadKernelChannel_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(11) & loadKernelChannel_CP_1349_elements(34) & loadKernelChannel_CP_1349_elements(44) & loadKernelChannel_CP_1349_elements(51) & loadKernelChannel_CP_1349_elements(58);
      gj_loadKernelChannel_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	64 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_sample_completed__ps
      -- CP-element group 16: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/aggregated_phi_sample_ack
      -- 
    -- Element group loadKernelChannel_CP_1349_elements(16) is bound as output of CP function.
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17: 	34 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	56 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (16) 
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_resize_1/index_resize_req
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_scale_1/$exit
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_scale_1/$entry
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/aggregated_phi_update_ack
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Sample/req
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_scale_1/scale_rename_ack
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_resized_1
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_scaled_1
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_computed_1
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_update_completed__ps
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_resize_1/$entry
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_scale_1/scale_rename_req
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_resize_1/$exit
      -- CP-element group 17: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_index_resize_1/index_resize_ack
      -- 
    req_1474_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1474_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(17), ack => array_obj_ref_468_index_offset_req_0); -- 
    -- Element group loadKernelChannel_CP_1349_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	9 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_loopback_trigger
      -- 
    loadKernelChannel_CP_1349_elements(18) <= loadKernelChannel_CP_1349_elements(9);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_loopback_sample_req
      -- CP-element group 19: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_loopback_sample_req_ps
      -- 
    phi_stmt_453_loopback_sample_req_1405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_loopback_sample_req_1405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(19), ack => phi_stmt_453_req_0); -- 
    -- Element group loadKernelChannel_CP_1349_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	10 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_entry_trigger
      -- 
    loadKernelChannel_CP_1349_elements(20) <= loadKernelChannel_CP_1349_elements(10);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_entry_sample_req
      -- CP-element group 21: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_entry_sample_req_ps
      -- 
    phi_stmt_453_entry_sample_req_1408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_453_entry_sample_req_1408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(21), ack => phi_stmt_453_req_1); -- 
    -- Element group loadKernelChannel_CP_1349_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_phi_mux_ack
      -- CP-element group 22: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/phi_stmt_453_phi_mux_ack_ps
      -- 
    phi_stmt_453_phi_mux_ack_1411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_453_ack_0, ack => loadKernelChannel_CP_1349_elements(22)); -- 
    -- CP-element group 23:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	25 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Sample/req
      -- CP-element group 23: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_sample_start__ps
      -- 
    req_1424_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1424_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(23), ack => nmycount_462_455_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1349_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_update_start__ps
      -- CP-element group 24: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_update_start_
      -- CP-element group 24: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Update/$entry
      -- CP-element group 24: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Update/req
      -- 
    req_1429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(24), ack => nmycount_462_455_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1349_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	23 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Sample/ack
      -- CP-element group 25: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_sample_completed__ps
      -- 
    ack_1425_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_462_455_buf_ack_0, ack => loadKernelChannel_CP_1349_elements(25)); -- 
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_update_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_nmycount_455_Update/ack
      -- 
    ack_1430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmycount_462_455_buf_ack_1, ack => loadKernelChannel_CP_1349_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Sample/req
      -- CP-element group 27: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Sample/$entry
      -- 
    req_1442_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1442_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(27), ack => start_add_456_buf_req_0); -- 
    -- Element group loadKernelChannel_CP_1349_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Update/$entry
      -- CP-element group 28: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Update/req
      -- CP-element group 28: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_update_start_
      -- 
    req_1447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(28), ack => start_add_456_buf_req_1); -- 
    -- Element group loadKernelChannel_CP_1349_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_sample_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Sample/$exit
      -- 
    ack_1443_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_456_buf_ack_0, ack => loadKernelChannel_CP_1349_elements(29)); -- 
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_update_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/R_start_add_456_update_completed_
      -- 
    ack_1448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => start_add_456_buf_ack_1, ack => loadKernelChannel_CP_1349_elements(30)); -- 
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	35 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	36 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_request/req
      -- CP-element group 31: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_request/$entry
      -- 
    req_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(31), ack => addr_of_469_final_reg_req_0); -- 
    loadKernelChannel_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(35) & loadKernelChannel_CP_1349_elements(36);
      gj_loadKernelChannel_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	11 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	40 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	37 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_complete/req
      -- CP-element group 32: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_update_start_
      -- CP-element group 32: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_complete/$entry
      -- 
    req_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(32), ack => addr_of_469_final_reg_req_1); -- 
    loadKernelChannel_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(11) & loadKernelChannel_CP_1349_elements(40);
      gj_loadKernelChannel_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_update_start
      -- CP-element group 33: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Update/req
      -- 
    req_1479_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1479_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(33), ack => array_obj_ref_468_index_offset_req_1); -- 
    loadKernelChannel_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(11) & loadKernelChannel_CP_1349_elements(36);
      gj_loadKernelChannel_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	17 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	64 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	15 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_sample_complete
      -- CP-element group 34: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Sample/ack
      -- 
    ack_1475_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_468_index_offset_ack_0, ack => loadKernelChannel_CP_1349_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	31 
    -- CP-element group 35:  members (8) 
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_final_index_sum_regn_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_root_address_calculated
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_offset_calculated
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_base_plus_offset/$entry
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_base_plus_offset/$exit
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_base_plus_offset/sum_rename_req
      -- CP-element group 35: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/array_obj_ref_468_base_plus_offset/sum_rename_ack
      -- 
    ack_1480_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_468_index_offset_ack_1, ack => loadKernelChannel_CP_1349_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	31 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_request/ack
      -- CP-element group 36: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_request/$exit
      -- 
    ack_1490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_469_final_reg_ack_0, ack => loadKernelChannel_CP_1349_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	32 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (19) 
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_addr_resize/$exit
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_complete/ack
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/addr_of_469_complete/$exit
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_addr_resize/base_resize_req
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_word_addrgen/root_register_req
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_word_addrgen/$entry
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_word_addrgen/root_register_ack
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_addr_resize/base_resize_ack
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_root_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_word_addrgen/$exit
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_address_resized
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_plus_offset/$entry
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_plus_offset/$exit
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_word_address_calculated
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_addr_resize/$entry
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_plus_offset/sum_rename_ack
      -- CP-element group 37: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_base_plus_offset/sum_rename_req
      -- 
    ack_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_469_final_reg_ack_1, ack => loadKernelChannel_CP_1349_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (5) 
      -- CP-element group 38: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/word_0/rr
      -- CP-element group 38: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/$entry
      -- CP-element group 38: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/word_0/$entry
      -- 
    rr_1528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(38), ack => ptr_deref_473_load_0_req_0); -- 
    loadKernelChannel_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(37) & loadKernelChannel_CP_1349_elements(40);
      gj_loadKernelChannel_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	47 
    -- CP-element group 39: 	54 
    -- CP-element group 39: 	61 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (5) 
      -- CP-element group 39: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/$entry
      -- CP-element group 39: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_update_start_
      -- CP-element group 39: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/word_0/$entry
      -- CP-element group 39: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/word_0/cr
      -- 
    cr_1539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(39), ack => ptr_deref_473_load_0_req_1); -- 
    loadKernelChannel_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(47) & loadKernelChannel_CP_1349_elements(54) & loadKernelChannel_CP_1349_elements(61);
      gj_loadKernelChannel_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	32 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (5) 
      -- CP-element group 40: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/word_0/$exit
      -- CP-element group 40: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/word_0/ra
      -- CP-element group 40: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Sample/word_access_start/$exit
      -- 
    ra_1529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_473_load_0_ack_0, ack => loadKernelChannel_CP_1349_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	46 
    -- CP-element group 41: 	53 
    -- CP-element group 41: 	60 
    -- CP-element group 41:  members (9) 
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/$exit
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/ptr_deref_473_Merge/merge_req
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/ptr_deref_473_Merge/merge_ack
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/word_0/$exit
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/word_access_complete/word_0/ca
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/ptr_deref_473_Merge/$entry
      -- CP-element group 41: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/ptr_deref_473_Update/ptr_deref_473_Merge/$exit
      -- 
    ca_1540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_473_load_0_ack_1, ack => loadKernelChannel_CP_1349_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Sample/req
      -- CP-element group 42: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_sample_start_
      -- 
    req_1553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(42), ack => W_send_to_1_481_delayed_13_0_493_inst_req_0); -- 
    loadKernelChannel_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(17) & loadKernelChannel_CP_1349_elements(44);
      gj_loadKernelChannel_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	47 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Update/req
      -- CP-element group 43: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_update_start_
      -- 
    req_1558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(43), ack => W_send_to_1_481_delayed_13_0_493_inst_req_1); -- 
    loadKernelChannel_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadKernelChannel_CP_1349_elements(47);
      gj_loadKernelChannel_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	15 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Sample/ack
      -- CP-element group 44: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_sample_completed_
      -- 
    ack_1554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_1_481_delayed_13_0_493_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_Update/ack
      -- CP-element group 45: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_495_update_completed_
      -- 
    ack_1559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_1_481_delayed_13_0_493_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	41 
    -- CP-element group 46: 	45 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Sample/$entry
      -- 
    req_1567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(46), ack => WPIPE_kernel_pipe1_497_inst_req_0); -- 
    loadKernelChannel_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(41) & loadKernelChannel_CP_1349_elements(45) & loadKernelChannel_CP_1349_elements(48);
      gj_loadKernelChannel_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	39 
    -- CP-element group 47: 	43 
    -- CP-element group 47:  members (6) 
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_update_start_
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Update/req
      -- CP-element group 47: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Sample/$exit
      -- 
    ack_1568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_497_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(47)); -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(47), ack => WPIPE_kernel_pipe1_497_inst_req_1); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	64 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe1_497_Update/ack
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe1_497_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	17 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Sample/req
      -- 
    req_1581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(49), ack => W_send_to_2_485_delayed_13_0_500_inst_req_0); -- 
    loadKernelChannel_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(17) & loadKernelChannel_CP_1349_elements(51);
      gj_loadKernelChannel_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	54 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Update/req
      -- CP-element group 50: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_update_start_
      -- CP-element group 50: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Update/$entry
      -- 
    req_1586_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1586_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(50), ack => W_send_to_2_485_delayed_13_0_500_inst_req_1); -- 
    loadKernelChannel_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadKernelChannel_CP_1349_elements(54);
      gj_loadKernelChannel_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	15 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Sample/$exit
      -- 
    ack_1582_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_2_485_delayed_13_0_500_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(51)); -- 
    -- CP-element group 52:  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_502_Update/ack
      -- 
    ack_1587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_2_485_delayed_13_0_500_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	41 
    -- CP-element group 53: 	52 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Sample/req
      -- CP-element group 53: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_sample_start_
      -- 
    req_1595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(53), ack => WPIPE_kernel_pipe2_504_inst_req_0); -- 
    loadKernelChannel_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(41) & loadKernelChannel_CP_1349_elements(52) & loadKernelChannel_CP_1349_elements(55);
      gj_loadKernelChannel_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	39 
    -- CP-element group 54: 	50 
    -- CP-element group 54:  members (6) 
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_update_start_
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Sample/ack
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Update/req
      -- 
    ack_1596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_504_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(54)); -- 
    req_1600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(54), ack => WPIPE_kernel_pipe2_504_inst_req_1); -- 
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	64 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe2_504_Update/$exit
      -- 
    ack_1601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe2_504_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	17 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_sample_start_
      -- CP-element group 56: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Sample/req
      -- 
    req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(56), ack => W_send_to_3_489_delayed_13_0_507_inst_req_0); -- 
    loadKernelChannel_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(17) & loadKernelChannel_CP_1349_elements(58);
      gj_loadKernelChannel_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	61 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_update_start_
      -- CP-element group 57: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Update/req
      -- CP-element group 57: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Update/$entry
      -- 
    req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1614_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(57), ack => W_send_to_3_489_delayed_13_0_507_inst_req_1); -- 
    loadKernelChannel_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadKernelChannel_CP_1349_elements(61);
      gj_loadKernelChannel_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	15 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Sample/ack
      -- 
    ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_3_489_delayed_13_0_507_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/assign_stmt_509_Update/$exit
      -- 
    ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_to_3_489_delayed_13_0_507_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	41 
    -- CP-element group 60: 	59 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Sample/req
      -- 
    req_1623_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1623_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(60), ack => WPIPE_kernel_pipe3_511_inst_req_0); -- 
    loadKernelChannel_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(41) & loadKernelChannel_CP_1349_elements(59) & loadKernelChannel_CP_1349_elements(62);
      gj_loadKernelChannel_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	62 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	39 
    -- CP-element group 61: 	57 
    -- CP-element group 61:  members (6) 
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_update_start_
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Sample/ack
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Update/req
      -- 
    ack_1624_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_511_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(61)); -- 
    req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1628_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(61), ack => WPIPE_kernel_pipe3_511_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	61 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/WPIPE_kernel_pipe3_511_Update/ack
      -- 
    ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_kernel_pipe3_511_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(62)); -- 
    -- CP-element group 63:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	11 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	12 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group loadKernelChannel_CP_1349_elements(63) is a control-delay.
    cp_element_63_delay: control_delay_element  generic map(name => " 63_delay", delay_value => 1)  port map(req => loadKernelChannel_CP_1349_elements(11), ack => loadKernelChannel_CP_1349_elements(63), clk => clk, reset =>reset);
    -- CP-element group 64:  join  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	16 
    -- CP-element group 64: 	34 
    -- CP-element group 64: 	48 
    -- CP-element group 64: 	55 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	8 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_450/do_while_stmt_451/do_while_stmt_451_loop_body/$exit
      -- 
    loadKernelChannel_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 37) := "loadKernelChannel_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= loadKernelChannel_CP_1349_elements(16) & loadKernelChannel_CP_1349_elements(34) & loadKernelChannel_CP_1349_elements(48) & loadKernelChannel_CP_1349_elements(55) & loadKernelChannel_CP_1349_elements(62);
      gj_loadKernelChannel_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	7 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_450/do_while_stmt_451/loop_exit/$exit
      -- CP-element group 65: 	 branch_block_stmt_450/do_while_stmt_451/loop_exit/ack
      -- 
    ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_451_branch_ack_0, ack => loadKernelChannel_CP_1349_elements(65)); -- 
    -- CP-element group 66:  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	7 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_450/do_while_stmt_451/loop_taken/$exit
      -- CP-element group 66: 	 branch_block_stmt_450/do_while_stmt_451/loop_taken/ack
      -- 
    ack_1638_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_451_branch_ack_1, ack => loadKernelChannel_CP_1349_elements(66)); -- 
    -- CP-element group 67:  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	5 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	3 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_450/do_while_stmt_451/$exit
      -- 
    loadKernelChannel_CP_1349_elements(67) <= loadKernelChannel_CP_1349_elements(5);
    -- CP-element group 68:  transition  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	3 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_sample_completed_
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_update_start_
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_Sample/$exit
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_Sample/ack
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_Update/$entry
      -- CP-element group 68: 	 assign_stmt_523/WPIPE_size_pipe_521_Update/req
      -- 
    ack_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_521_inst_ack_0, ack => loadKernelChannel_CP_1349_elements(68)); -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadKernelChannel_CP_1349_elements(68), ack => WPIPE_size_pipe_521_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (5) 
      -- CP-element group 69: 	 $exit
      -- CP-element group 69: 	 assign_stmt_523/$exit
      -- CP-element group 69: 	 assign_stmt_523/WPIPE_size_pipe_521_update_completed_
      -- CP-element group 69: 	 assign_stmt_523/WPIPE_size_pipe_521_Update/$exit
      -- CP-element group 69: 	 assign_stmt_523/WPIPE_size_pipe_521_Update/ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_size_pipe_521_inst_ack_1, ack => loadKernelChannel_CP_1349_elements(69)); -- 
    loadKernelChannel_do_while_stmt_451_terminator_1639: loop_terminator -- 
      generic map (name => " loadKernelChannel_do_while_stmt_451_terminator_1639", max_iterations_in_flight =>15) 
      port map(loop_body_exit => loadKernelChannel_CP_1349_elements(8),loop_continue => loadKernelChannel_CP_1349_elements(66),loop_terminate => loadKernelChannel_CP_1349_elements(65),loop_back => loadKernelChannel_CP_1349_elements(6),loop_exit => loadKernelChannel_CP_1349_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_453_phi_seq_1449_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= loadKernelChannel_CP_1349_elements(18);
      loadKernelChannel_CP_1349_elements(23)<= src_sample_reqs(0);
      src_sample_acks(0)  <= loadKernelChannel_CP_1349_elements(25);
      loadKernelChannel_CP_1349_elements(24)<= src_update_reqs(0);
      src_update_acks(0)  <= loadKernelChannel_CP_1349_elements(26);
      loadKernelChannel_CP_1349_elements(19) <= phi_mux_reqs(0);
      triggers(1)  <= loadKernelChannel_CP_1349_elements(20);
      loadKernelChannel_CP_1349_elements(27)<= src_sample_reqs(1);
      src_sample_acks(1)  <= loadKernelChannel_CP_1349_elements(29);
      loadKernelChannel_CP_1349_elements(28)<= src_update_reqs(1);
      src_update_acks(1)  <= loadKernelChannel_CP_1349_elements(30);
      loadKernelChannel_CP_1349_elements(21) <= phi_mux_reqs(1);
      phi_stmt_453_phi_seq_1449 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_453_phi_seq_1449") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => loadKernelChannel_CP_1349_elements(13), 
          phi_sample_ack => loadKernelChannel_CP_1349_elements(16), 
          phi_update_req => loadKernelChannel_CP_1349_elements(15), 
          phi_update_ack => loadKernelChannel_CP_1349_elements(17), 
          phi_mux_ack => loadKernelChannel_CP_1349_elements(22), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1391_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= loadKernelChannel_CP_1349_elements(9);
        preds(1)  <= loadKernelChannel_CP_1349_elements(10);
        entry_tmerge_1391 : transition_merge -- 
          generic map(name => " entry_tmerge_1391")
          port map (preds => preds, symbol_out => loadKernelChannel_CP_1349_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u1_u1_482_wire : std_logic_vector(0 downto 0);
    signal SHL_u16_u16_418_wire : std_logic_vector(15 downto 0);
    signal SHL_u16_u16_431_wire : std_logic_vector(15 downto 0);
    signal SUB_u32_u32_518_wire : std_logic_vector(31 downto 0);
    signal ULT_u32_u1_485_wire : std_logic_vector(0 downto 0);
    signal ULT_u32_u1_519_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_468_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_468_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_468_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_468_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_468_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_468_root_address : std_logic_vector(13 downto 0);
    signal ea1_426 : std_logic_vector(31 downto 0);
    signal ea2_434 : std_logic_vector(31 downto 0);
    signal ea3_440 : std_logic_vector(31 downto 0);
    signal fetch_addr_470 : std_logic_vector(31 downto 0);
    signal first_fill_445 : std_logic_vector(0 downto 0);
    signal konst_417_wire_constant : std_logic_vector(15 downto 0);
    signal konst_430_wire_constant : std_logic_vector(15 downto 0);
    signal konst_443_wire_constant : std_logic_vector(31 downto 0);
    signal konst_460_wire_constant : std_logic_vector(31 downto 0);
    signal konst_517_wire_constant : std_logic_vector(31 downto 0);
    signal my_fetch_474 : std_logic_vector(63 downto 0);
    signal mycount_453 : std_logic_vector(31 downto 0);
    signal nmycount_462 : std_logic_vector(31 downto 0);
    signal nmycount_462_455_buffered : std_logic_vector(31 downto 0);
    signal ptr_deref_473_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_473_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_473_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_473_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_473_word_offset_0 : std_logic_vector(13 downto 0);
    signal row_size_420 : std_logic_vector(15 downto 0);
    signal send_to_1_479 : std_logic_vector(0 downto 0);
    signal send_to_1_481_delayed_13_0_495 : std_logic_vector(0 downto 0);
    signal send_to_2_485_delayed_13_0_502 : std_logic_vector(0 downto 0);
    signal send_to_2_487 : std_logic_vector(0 downto 0);
    signal send_to_3_489_delayed_13_0_509 : std_logic_vector(0 downto 0);
    signal send_to_3_492 : std_logic_vector(0 downto 0);
    signal start_add_456_buffered : std_logic_vector(31 downto 0);
    signal start_next_449 : std_logic_vector(7 downto 0);
    signal type_cast_424_wire : std_logic_vector(31 downto 0);
    signal type_cast_432_wire : std_logic_vector(31 downto 0);
    signal type_cast_438_wire : std_logic_vector(31 downto 0);
    signal type_cast_467_resized : std_logic_vector(13 downto 0);
    signal type_cast_467_scaled : std_logic_vector(13 downto 0);
    signal type_cast_467_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_468_constant_part_of_offset <= "00000000000000";
    array_obj_ref_468_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_468_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_468_resized_base_address <= "00000000000000";
    konst_417_wire_constant <= "0000000000000001";
    konst_430_wire_constant <= "0000000000000001";
    konst_443_wire_constant <= "00000000000000000000000000000000";
    konst_460_wire_constant <= "00000000000000000000000000000001";
    konst_517_wire_constant <= "00000000000000000000000000000001";
    ptr_deref_473_word_offset_0 <= "00000000000000";
    phi_stmt_453: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nmycount_462_455_buffered & start_add_456_buffered;
      req <= phi_stmt_453_req_0 & phi_stmt_453_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_453",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_453_ack_0,
          idata => idata,
          odata => mycount_453,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_453
    W_send_to_1_481_delayed_13_0_493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_to_1_481_delayed_13_0_493_inst_req_0;
      W_send_to_1_481_delayed_13_0_493_inst_ack_0<= wack(0);
      rreq(0) <= W_send_to_1_481_delayed_13_0_493_inst_req_1;
      W_send_to_1_481_delayed_13_0_493_inst_ack_1<= rack(0);
      W_send_to_1_481_delayed_13_0_493_inst : InterlockBuffer generic map ( -- 
        name => "W_send_to_1_481_delayed_13_0_493_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_to_1_479,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_to_1_481_delayed_13_0_495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_to_2_485_delayed_13_0_500_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_to_2_485_delayed_13_0_500_inst_req_0;
      W_send_to_2_485_delayed_13_0_500_inst_ack_0<= wack(0);
      rreq(0) <= W_send_to_2_485_delayed_13_0_500_inst_req_1;
      W_send_to_2_485_delayed_13_0_500_inst_ack_1<= rack(0);
      W_send_to_2_485_delayed_13_0_500_inst : InterlockBuffer generic map ( -- 
        name => "W_send_to_2_485_delayed_13_0_500_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_to_2_487,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_to_2_485_delayed_13_0_502,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_to_3_489_delayed_13_0_507_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_to_3_489_delayed_13_0_507_inst_req_0;
      W_send_to_3_489_delayed_13_0_507_inst_ack_0<= wack(0);
      rreq(0) <= W_send_to_3_489_delayed_13_0_507_inst_req_1;
      W_send_to_3_489_delayed_13_0_507_inst_ack_1<= rack(0);
      W_send_to_3_489_delayed_13_0_507_inst : InterlockBuffer generic map ( -- 
        name => "W_send_to_3_489_delayed_13_0_507_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_to_3_492,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_to_3_489_delayed_13_0_509,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_469_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_469_final_reg_req_0;
      addr_of_469_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_469_final_reg_req_1;
      addr_of_469_final_reg_ack_1<= rack(0);
      addr_of_469_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_469_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_468_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmycount_462_455_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmycount_462_455_buf_req_0;
      nmycount_462_455_buf_ack_0<= wack(0);
      rreq(0) <= nmycount_462_455_buf_req_1;
      nmycount_462_455_buf_ack_1<= rack(0);
      nmycount_462_455_buf : InterlockBuffer generic map ( -- 
        name => "nmycount_462_455_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmycount_462,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmycount_462_455_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    start_add_456_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= start_add_456_buf_req_0;
      start_add_456_buf_ack_0<= wack(0);
      rreq(0) <= start_add_456_buf_req_1;
      start_add_456_buf_ack_1<= rack(0);
      start_add_456_buf : InterlockBuffer generic map ( -- 
        name => "start_add_456_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => start_add_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => start_add_456_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_424_inst
    process(row_size_420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_420(15 downto 0);
      type_cast_424_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_432_inst
    process(SHL_u16_u16_431_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := SHL_u16_u16_431_wire(15 downto 0);
      type_cast_432_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_438_inst
    process(row_size_420) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := row_size_420(15 downto 0);
      type_cast_438_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_467_inst
    process(mycount_453) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := mycount_453(31 downto 0);
      type_cast_467_wire <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_468_index_1_rename
    process(type_cast_467_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_467_resized;
      ov(13 downto 0) := iv;
      type_cast_467_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_468_index_1_resize
    process(type_cast_467_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_467_wire;
      ov := iv(13 downto 0);
      type_cast_467_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_468_root_address_inst
    process(array_obj_ref_468_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_468_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_468_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_473_addr_0
    process(ptr_deref_473_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_473_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_473_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_473_base_resize
    process(fetch_addr_470) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr_470;
      ov := iv(13 downto 0);
      ptr_deref_473_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_473_gather_scatter
    process(ptr_deref_473_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_473_data_0;
      ov(63 downto 0) := iv;
      my_fetch_474 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_473_root_address_inst
    process(ptr_deref_473_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_473_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_473_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_451_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u32_u1_519_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_451_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_451_branch_req_0,
          ack0 => do_while_stmt_451_branch_ack_0,
          ack1 => do_while_stmt_451_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_419_inst
    process(num_chl_buffer, SHL_u16_u16_418_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(num_chl_buffer, SHL_u16_u16_418_wire, tmp_var);
      row_size_420 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_425_inst
    process(start_add_buffer, type_cast_424_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_424_wire, tmp_var);
      ea1_426 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_433_inst
    process(start_add_buffer, type_cast_432_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(start_add_buffer, type_cast_432_wire, tmp_var);
      ea2_434 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_439_inst
    process(ea2_434, type_cast_438_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ea2_434, type_cast_438_wire, tmp_var);
      ea3_440 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_461_inst
    process(mycount_453) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mycount_453, konst_460_wire_constant, tmp_var);
      nmycount_462 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_486_inst
    process(NOT_u1_u1_482_wire, ULT_u32_u1_485_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_482_wire, ULT_u32_u1_485_wire, tmp_var);
      send_to_2_487 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_444_inst
    process(start_add_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(start_add_buffer, konst_443_wire_constant, tmp_var);
      first_fill_445 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_482_inst
    process(send_to_1_479) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", send_to_1_479, tmp_var);
      NOT_u1_u1_482_wire <= tmp_var; -- 
    end process;
    -- binary operator SHL_u16_u16_418_inst
    process(num_chl_buffer) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(num_chl_buffer, konst_417_wire_constant, tmp_var);
      SHL_u16_u16_418_wire <= tmp_var; --
    end process;
    -- binary operator SHL_u16_u16_431_inst
    process(row_size_420) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntSHL_proc(row_size_420, konst_430_wire_constant, tmp_var);
      SHL_u16_u16_431_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_518_inst
    process(ea3_440) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(ea3_440, konst_517_wire_constant, tmp_var);
      SUB_u32_u32_518_wire <= tmp_var; --
    end process;
    -- binary operator UGE_u32_u1_491_inst
    process(mycount_453, ea2_434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(mycount_453, ea2_434, tmp_var);
      send_to_3_492 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_478_inst
    process(mycount_453, ea1_426) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_453, ea1_426, tmp_var);
      send_to_1_479 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_485_inst
    process(mycount_453, ea2_434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_453, ea2_434, tmp_var);
      ULT_u32_u1_485_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_519_inst
    process(mycount_453, SUB_u32_u32_518_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(mycount_453, SUB_u32_u32_518_wire, tmp_var);
      ULT_u32_u1_519_wire <= tmp_var; --
    end process;
    -- shared split operator group (15) : array_obj_ref_468_index_offset 
    ApIntAdd_group_15: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_467_scaled;
      array_obj_ref_468_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_468_index_offset_req_0;
      array_obj_ref_468_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_468_index_offset_req_1;
      array_obj_ref_468_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_15_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_15_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_15",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared load operator group (0) : ptr_deref_473_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 6);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_473_load_0_req_0;
      ptr_deref_473_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_473_load_0_req_1;
      ptr_deref_473_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_473_word_address_0;
      ptr_deref_473_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(13 downto 0),
          mtag => memory_space_1_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(63 downto 0),
          mtag => memory_space_1_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_input_done_pipe_448_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_input_done_pipe_448_inst_req_0;
      RPIPE_input_done_pipe_448_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_input_done_pipe_448_inst_req_1;
      RPIPE_input_done_pipe_448_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not first_fill_445(0);
      start_next_449 <= data_out(7 downto 0);
      input_done_pipe_read_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_read_0: InputPortRevised -- 
        generic map ( name => "input_done_pipe_read_0", data_width => 8,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => input_done_pipe_pipe_read_req(0),
          oack => input_done_pipe_pipe_read_ack(0),
          odata => input_done_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_kernel_pipe1_497_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe1_497_inst_req_0;
      WPIPE_kernel_pipe1_497_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe1_497_inst_req_1;
      WPIPE_kernel_pipe1_497_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_1_481_delayed_13_0_495(0);
      data_in <= my_fetch_474;
      kernel_pipe1_write_0_gI: SplitGuardInterface generic map(name => "kernel_pipe1_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe1_write_0: OutputPortRevised -- 
        generic map ( name => "kernel_pipe1", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe1_pipe_write_req(0),
          oack => kernel_pipe1_pipe_write_ack(0),
          odata => kernel_pipe1_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_kernel_pipe2_504_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe2_504_inst_req_0;
      WPIPE_kernel_pipe2_504_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe2_504_inst_req_1;
      WPIPE_kernel_pipe2_504_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_2_485_delayed_13_0_502(0);
      data_in <= my_fetch_474;
      kernel_pipe2_write_1_gI: SplitGuardInterface generic map(name => "kernel_pipe2_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe2_write_1: OutputPortRevised -- 
        generic map ( name => "kernel_pipe2", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe2_pipe_write_req(0),
          oack => kernel_pipe2_pipe_write_ack(0),
          odata => kernel_pipe2_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_kernel_pipe3_511_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_kernel_pipe3_511_inst_req_0;
      WPIPE_kernel_pipe3_511_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_kernel_pipe3_511_inst_req_1;
      WPIPE_kernel_pipe3_511_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_to_3_489_delayed_13_0_509(0);
      data_in <= my_fetch_474;
      kernel_pipe3_write_2_gI: SplitGuardInterface generic map(name => "kernel_pipe3_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      kernel_pipe3_write_2: OutputPortRevised -- 
        generic map ( name => "kernel_pipe3", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => kernel_pipe3_pipe_write_req(0),
          oack => kernel_pipe3_pipe_write_ack(0),
          odata => kernel_pipe3_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_size_pipe_521_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_size_pipe_521_inst_req_0;
      WPIPE_size_pipe_521_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_size_pipe_521_inst_req_1;
      WPIPE_size_pipe_521_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= num_chl_buffer;
      size_pipe_write_3_gI: SplitGuardInterface generic map(name => "size_pipe_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      size_pipe_write_3: OutputPortRevised -- 
        generic map ( name => "size_pipe", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => size_pipe_pipe_write_req(0),
          oack => size_pipe_pipe_write_ack(0),
          odata => size_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end loadKernelChannel_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendB is -- 
  generic (tag_length : integer); 
  port ( -- 
    size : in  std_logic_vector(31 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendB;
architecture sendB_arch of sendB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal size_buffer :  std_logic_vector(31 downto 0);
  signal size_update_enable: Boolean;
  -- output port buffer signals
  signal sendB_CP_1657_start: Boolean;
  signal sendB_CP_1657_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_609_inst_req_1 : boolean;
  signal type_cast_599_inst_req_1 : boolean;
  signal ptr_deref_595_load_0_req_1 : boolean;
  signal if_stmt_534_branch_ack_0 : boolean;
  signal ptr_deref_595_load_0_ack_1 : boolean;
  signal type_cast_599_inst_ack_0 : boolean;
  signal type_cast_649_inst_req_1 : boolean;
  signal type_cast_561_inst_ack_1 : boolean;
  signal type_cast_609_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_1 : boolean;
  signal array_obj_ref_590_index_offset_ack_0 : boolean;
  signal type_cast_669_inst_req_0 : boolean;
  signal array_obj_ref_590_index_offset_req_0 : boolean;
  signal array_obj_ref_590_index_offset_ack_1 : boolean;
  signal addr_of_591_final_reg_ack_1 : boolean;
  signal type_cast_669_inst_ack_0 : boolean;
  signal type_cast_599_inst_req_0 : boolean;
  signal if_stmt_534_branch_ack_1 : boolean;
  signal type_cast_561_inst_ack_0 : boolean;
  signal type_cast_609_inst_req_0 : boolean;
  signal ptr_deref_595_load_0_req_0 : boolean;
  signal type_cast_649_inst_ack_0 : boolean;
  signal type_cast_669_inst_ack_1 : boolean;
  signal array_obj_ref_590_index_offset_req_1 : boolean;
  signal type_cast_629_inst_req_1 : boolean;
  signal type_cast_619_inst_ack_1 : boolean;
  signal type_cast_619_inst_req_1 : boolean;
  signal type_cast_649_inst_req_0 : boolean;
  signal type_cast_639_inst_ack_0 : boolean;
  signal type_cast_629_inst_ack_1 : boolean;
  signal type_cast_609_inst_ack_0 : boolean;
  signal type_cast_599_inst_ack_1 : boolean;
  signal addr_of_591_final_reg_req_1 : boolean;
  signal ptr_deref_595_load_0_ack_0 : boolean;
  signal type_cast_659_inst_ack_1 : boolean;
  signal type_cast_561_inst_req_0 : boolean;
  signal type_cast_659_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_683_inst_ack_1 : boolean;
  signal type_cast_649_inst_ack_1 : boolean;
  signal type_cast_659_inst_ack_0 : boolean;
  signal type_cast_619_inst_ack_0 : boolean;
  signal addr_of_591_final_reg_ack_0 : boolean;
  signal type_cast_629_inst_ack_0 : boolean;
  signal type_cast_639_inst_ack_1 : boolean;
  signal type_cast_639_inst_req_1 : boolean;
  signal type_cast_639_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_692_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_692_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_692_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_692_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_674_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_674_inst_req_1 : boolean;
  signal type_cast_659_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_671_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_671_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_677_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_671_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_677_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_674_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_671_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_674_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_683_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_677_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_689_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_689_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_683_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_683_inst_req_1 : boolean;
  signal if_stmt_706_branch_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_677_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_686_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_686_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_680_inst_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_680_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_680_inst_req_0 : boolean;
  signal type_cast_629_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_680_inst_req_1 : boolean;
  signal if_stmt_706_branch_ack_1 : boolean;
  signal if_stmt_706_branch_ack_0 : boolean;
  signal WPIPE_maxpool_output_pipe_686_inst_req_1 : boolean;
  signal WPIPE_maxpool_output_pipe_686_inst_ack_1 : boolean;
  signal WPIPE_maxpool_output_pipe_689_inst_req_0 : boolean;
  signal WPIPE_maxpool_output_pipe_689_inst_ack_0 : boolean;
  signal type_cast_619_inst_req_0 : boolean;
  signal phi_stmt_578_req_0 : boolean;
  signal type_cast_669_inst_req_1 : boolean;
  signal if_stmt_534_branch_req_0 : boolean;
  signal type_cast_584_inst_req_0 : boolean;
  signal type_cast_584_inst_ack_0 : boolean;
  signal type_cast_584_inst_req_1 : boolean;
  signal type_cast_584_inst_ack_1 : boolean;
  signal phi_stmt_578_req_1 : boolean;
  signal phi_stmt_578_ack_0 : boolean;
  signal addr_of_591_final_reg_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= size;
  size_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendB_CP_1657_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1657_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendB_CP_1657_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendB_CP_1657_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendB_CP_1657: Block -- control-path 
    signal sendB_CP_1657_elements: BooleanArray(59 downto 0);
    -- 
  begin -- 
    sendB_CP_1657_elements(0) <= sendB_CP_1657_start;
    sendB_CP_1657_symbol <= sendB_CP_1657_elements(59);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (15) 
      -- CP-element group 0: 	 branch_block_stmt_527/assign_stmt_533/$entry
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534__entry__
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_if_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_else_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_527/assign_stmt_533__entry__
      -- CP-element group 0: 	 branch_block_stmt_527/assign_stmt_533/$exit
      -- CP-element group 0: 	 branch_block_stmt_527/assign_stmt_533__exit__
      -- CP-element group 0: 	 branch_block_stmt_527/branch_block_stmt_527__entry__
      -- CP-element group 0: 	 branch_block_stmt_527/$entry
      -- CP-element group 0: 	 branch_block_stmt_527/R_cmp68_535_place
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_eval_test/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_527/if_stmt_534_eval_test/$entry
      -- 
    branch_req_1695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(0), ack => if_stmt_534_branch_req_0); -- 
    -- CP-element group 1:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (18) 
      -- CP-element group 1: 	 branch_block_stmt_527/merge_stmt_540__exit__
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575__entry__
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_527/if_stmt_534_if_link/if_choice_transition
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_527/if_stmt_534_if_link/$exit
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_update_start_
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/$entry
      -- CP-element group 1: 	 branch_block_stmt_527/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 1: 	 branch_block_stmt_527/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 1: 	 branch_block_stmt_527/entry_bbx_xnph
      -- CP-element group 1: 	 branch_block_stmt_527/merge_stmt_540_PhiReqMerge
      -- CP-element group 1: 	 branch_block_stmt_527/merge_stmt_540_PhiAck/$entry
      -- CP-element group 1: 	 branch_block_stmt_527/merge_stmt_540_PhiAck/$exit
      -- CP-element group 1: 	 branch_block_stmt_527/merge_stmt_540_PhiAck/dummy
      -- 
    if_choice_transition_1700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_534_branch_ack_1, ack => sendB_CP_1657_elements(1)); -- 
    cr_1722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(1), ack => type_cast_561_inst_req_1); -- 
    rr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1717_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(1), ack => type_cast_561_inst_req_0); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	59 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_527/if_stmt_534_else_link/else_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_527/if_stmt_534_else_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_527/entry_forx_xend
      -- CP-element group 2: 	 branch_block_stmt_527/entry_forx_xend_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_527/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_1704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_534_branch_ack_0, ack => sendB_CP_1657_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_sample_completed_
      -- 
    ra_1718_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_0, ack => sendB_CP_1657_elements(3)); -- 
    -- CP-element group 4:  transition  place  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	53 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_527/bbx_xnph_forx_xbody
      -- CP-element group 4: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575__exit__
      -- CP-element group 4: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_Update/ca
      -- CP-element group 4: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/type_cast_561_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_527/assign_stmt_546_to_assign_stmt_575/$exit
      -- CP-element group 4: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/$entry
      -- CP-element group 4: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/$entry
      -- 
    ca_1723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_561_inst_ack_1, ack => sendB_CP_1657_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	58 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	50 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_sample_complete
      -- CP-element group 5: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Sample/ack
      -- 
    ack_1752_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_590_index_offset_ack_0, ack => sendB_CP_1657_elements(5)); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	58 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_request/$entry
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_offset_calculated
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_base_plus_offset/$entry
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_base_plus_offset/sum_rename_ack
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_root_address_calculated
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_base_plus_offset/sum_rename_req
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_base_plus_offset/$exit
      -- CP-element group 6: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_request/req
      -- 
    ack_1757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_590_index_offset_ack_1, ack => sendB_CP_1657_elements(6)); -- 
    req_1766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(6), ack => addr_of_591_final_reg_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_request/$exit
      -- CP-element group 7: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_request/ack
      -- CP-element group 7: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_sample_completed_
      -- 
    ack_1767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_591_final_reg_ack_0, ack => sendB_CP_1657_elements(7)); -- 
    -- CP-element group 8:  join  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	58 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (24) 
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_word_addrgen/root_register_ack
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_plus_offset/sum_rename_ack
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_word_addrgen/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_plus_offset/sum_rename_req
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_word_addrgen/$exit
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_word_addrgen/root_register_req
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_complete/ack
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_addr_resize/base_resize_ack
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/word_0/rr
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_plus_offset/$exit
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_addr_resize/$exit
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_plus_offset/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_addr_resize/base_resize_req
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/word_0/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_addr_resize/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_address_resized
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/$entry
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_root_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_word_address_calculated
      -- CP-element group 8: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_base_address_calculated
      -- 
    ack_1772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_591_final_reg_ack_1, ack => sendB_CP_1657_elements(8)); -- 
    rr_1805_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1805_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(8), ack => ptr_deref_595_load_0_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Sample/$exit
      -- 
    ra_1806_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_load_0_ack_0, ack => sendB_CP_1657_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	58 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	17 
    -- CP-element group 10: 	19 
    -- CP-element group 10: 	21 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	25 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (33) 
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/ptr_deref_595_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/ptr_deref_595_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/ptr_deref_595_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Sample/rr
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/ptr_deref_595_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_update_completed_
      -- 
    ca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_load_0_ack_1, ack => sendB_CP_1657_elements(10)); -- 
    rr_1858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_619_inst_req_0); -- 
    rr_1872_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1872_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_629_inst_req_0); -- 
    rr_1886_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1886_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_639_inst_req_0); -- 
    rr_1900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_649_inst_req_0); -- 
    rr_1914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_659_inst_req_0); -- 
    rr_1928_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1928_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_669_inst_req_0); -- 
    rr_1844_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1844_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_609_inst_req_0); -- 
    rr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(10), ack => type_cast_599_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_sample_completed_
      -- 
    ra_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_0, ack => sendB_CP_1657_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	58 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	47 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_update_completed_
      -- 
    ca_1836_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_599_inst_ack_1, ack => sendB_CP_1657_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Sample/$exit
      -- 
    ra_1845_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_609_inst_ack_0, ack => sendB_CP_1657_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	44 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_update_completed_
      -- 
    ca_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_609_inst_ack_1, ack => sendB_CP_1657_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Sample/$exit
      -- 
    ra_1859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_619_inst_ack_0, ack => sendB_CP_1657_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	58 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Update/$exit
      -- 
    ca_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_619_inst_ack_1, ack => sendB_CP_1657_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	10 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Sample/ra
      -- 
    ra_1873_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_629_inst_ack_0, ack => sendB_CP_1657_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	58 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	38 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Update/$exit
      -- 
    ca_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_629_inst_ack_1, ack => sendB_CP_1657_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Sample/ra
      -- CP-element group 19: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Sample/$exit
      -- 
    ra_1887_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_0, ack => sendB_CP_1657_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	35 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Update/ca
      -- CP-element group 20: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Update/$exit
      -- 
    ca_1892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_639_inst_ack_1, ack => sendB_CP_1657_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_sample_completed_
      -- 
    ra_1901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_0, ack => sendB_CP_1657_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	58 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	32 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Update/ca
      -- 
    ca_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_649_inst_ack_1, ack => sendB_CP_1657_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Sample/ra
      -- 
    ra_1915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_0, ack => sendB_CP_1657_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	58 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Update/ca
      -- CP-element group 24: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Update/$exit
      -- 
    ca_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_659_inst_ack_1, ack => sendB_CP_1657_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	10 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Sample/ra
      -- CP-element group 25: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_sample_completed_
      -- 
    ra_1929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_0, ack => sendB_CP_1657_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	58 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Update/$exit
      -- 
    ca_1934_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_669_inst_ack_1, ack => sendB_CP_1657_elements(26)); -- 
    req_1942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(26), ack => WPIPE_maxpool_output_pipe_671_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Update/req
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_update_start_
      -- 
    ack_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_671_inst_ack_0, ack => sendB_CP_1657_elements(27)); -- 
    req_1947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(27), ack => WPIPE_maxpool_output_pipe_671_inst_req_1); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_671_Update/$exit
      -- 
    ack_1948_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_671_inst_ack_1, ack => sendB_CP_1657_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	24 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Sample/req
      -- 
    req_1956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(29), ack => WPIPE_maxpool_output_pipe_674_inst_req_0); -- 
    sendB_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(28) & sendB_CP_1657_elements(24);
      gj_sendB_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  output  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (6) 
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_update_start_
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Update/req
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Sample/ack
      -- 
    ack_1957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_674_inst_ack_0, ack => sendB_CP_1657_elements(30)); -- 
    req_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(30), ack => WPIPE_maxpool_output_pipe_674_inst_req_1); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Update/ack
      -- CP-element group 31: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_674_Update/$exit
      -- 
    ack_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_674_inst_ack_1, ack => sendB_CP_1657_elements(31)); -- 
    -- CP-element group 32:  join  transition  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: 	22 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Sample/req
      -- CP-element group 32: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Sample/$entry
      -- 
    req_1970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(32), ack => WPIPE_maxpool_output_pipe_677_inst_req_0); -- 
    sendB_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(31) & sendB_CP_1657_elements(22);
      gj_sendB_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	32 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_update_start_
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Update/req
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Sample/$exit
      -- 
    ack_1971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_677_inst_ack_0, ack => sendB_CP_1657_elements(33)); -- 
    req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(33), ack => WPIPE_maxpool_output_pipe_677_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_677_Update/$exit
      -- 
    ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_677_inst_ack_1, ack => sendB_CP_1657_elements(34)); -- 
    -- CP-element group 35:  join  transition  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	20 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Sample/req
      -- 
    req_1984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(35), ack => WPIPE_maxpool_output_pipe_680_inst_req_0); -- 
    sendB_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(20) & sendB_CP_1657_elements(34);
      gj_sendB_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Sample/ack
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_update_start_
      -- CP-element group 36: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Update/req
      -- 
    ack_1985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_680_inst_ack_0, ack => sendB_CP_1657_elements(36)); -- 
    req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1989_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(36), ack => WPIPE_maxpool_output_pipe_680_inst_req_1); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Update/ack
      -- CP-element group 37: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_680_Update/$exit
      -- 
    ack_1990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_680_inst_ack_1, ack => sendB_CP_1657_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	18 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Sample/req
      -- 
    req_1998_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1998_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(38), ack => WPIPE_maxpool_output_pipe_683_inst_req_0); -- 
    sendB_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(18) & sendB_CP_1657_elements(37);
      gj_sendB_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (6) 
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Update/req
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_update_start_
      -- CP-element group 39: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Sample/$exit
      -- 
    ack_1999_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_683_inst_ack_0, ack => sendB_CP_1657_elements(39)); -- 
    req_2003_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2003_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(39), ack => WPIPE_maxpool_output_pipe_683_inst_req_1); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_683_Update/$exit
      -- 
    ack_2004_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_683_inst_ack_1, ack => sendB_CP_1657_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Sample/req
      -- CP-element group 41: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Sample/$entry
      -- 
    req_2012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(41), ack => WPIPE_maxpool_output_pipe_686_inst_req_0); -- 
    sendB_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(16) & sendB_CP_1657_elements(40);
      gj_sendB_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (6) 
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_update_start_
      -- CP-element group 42: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Update/req
      -- 
    ack_2013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_686_inst_ack_0, ack => sendB_CP_1657_elements(42)); -- 
    req_2017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(42), ack => WPIPE_maxpool_output_pipe_686_inst_req_1); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_686_Update/ack
      -- 
    ack_2018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_686_inst_ack_1, ack => sendB_CP_1657_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	14 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Sample/req
      -- 
    req_2026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(44), ack => WPIPE_maxpool_output_pipe_689_inst_req_0); -- 
    sendB_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(14) & sendB_CP_1657_elements(43);
      gj_sendB_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_update_start_
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Update/req
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Sample/ack
      -- 
    ack_2027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_689_inst_ack_0, ack => sendB_CP_1657_elements(45)); -- 
    req_2031_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2031_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(45), ack => WPIPE_maxpool_output_pipe_689_inst_req_1); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Update/ack
      -- CP-element group 46: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_689_Update/$exit
      -- 
    ack_2032_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_689_inst_ack_1, ack => sendB_CP_1657_elements(46)); -- 
    -- CP-element group 47:  join  transition  output  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	12 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_sample_start_
      -- CP-element group 47: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Sample/req
      -- CP-element group 47: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Sample/$entry
      -- 
    req_2040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(47), ack => WPIPE_maxpool_output_pipe_692_inst_req_0); -- 
    sendB_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(12) & sendB_CP_1657_elements(46);
      gj_sendB_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (6) 
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Update/req
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_update_start_
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Sample/ack
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Update/$entry
      -- CP-element group 48: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_sample_completed_
      -- 
    ack_2041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_692_inst_ack_0, ack => sendB_CP_1657_elements(48)); -- 
    req_2045_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2045_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(48), ack => WPIPE_maxpool_output_pipe_692_inst_req_1); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Update/ack
      -- CP-element group 49: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/WPIPE_maxpool_output_pipe_692_Update/$exit
      -- 
    ack_2046_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_maxpool_output_pipe_692_inst_ack_1, ack => sendB_CP_1657_elements(49)); -- 
    -- CP-element group 50:  branch  join  transition  place  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	5 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (10) 
      -- CP-element group 50: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/$exit
      -- CP-element group 50: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705__exit__
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706__entry__
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_dead_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_eval_test/branch_req
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_eval_test/$entry
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_eval_test/$exit
      -- CP-element group 50: 	 branch_block_stmt_527/R_exitcond1_707_place
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_if_link/$entry
      -- CP-element group 50: 	 branch_block_stmt_527/if_stmt_706_else_link/$entry
      -- 
    branch_req_2054_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2054_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(50), ack => if_stmt_706_branch_req_0); -- 
    sendB_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(5) & sendB_CP_1657_elements(49);
      gj_sendB_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  merge  transition  place  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	59 
    -- CP-element group 51:  members (13) 
      -- CP-element group 51: 	 branch_block_stmt_527/merge_stmt_712__exit__
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xendx_xloopexit_forx_xend
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 51: 	 branch_block_stmt_527/if_stmt_706_if_link/$exit
      -- CP-element group 51: 	 branch_block_stmt_527/if_stmt_706_if_link/if_choice_transition
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 51: 	 branch_block_stmt_527/merge_stmt_712_PhiReqMerge
      -- CP-element group 51: 	 branch_block_stmt_527/merge_stmt_712_PhiAck/$entry
      -- CP-element group 51: 	 branch_block_stmt_527/merge_stmt_712_PhiAck/$exit
      -- CP-element group 51: 	 branch_block_stmt_527/merge_stmt_712_PhiAck/dummy
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 51: 	 branch_block_stmt_527/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_2059_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_706_branch_ack_1, ack => sendB_CP_1657_elements(51)); -- 
    -- CP-element group 52:  fork  transition  place  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: 	55 
    -- CP-element group 52:  members (12) 
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody
      -- CP-element group 52: 	 branch_block_stmt_527/if_stmt_706_else_link/else_choice_transition
      -- CP-element group 52: 	 branch_block_stmt_527/if_stmt_706_else_link/$exit
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Sample/rr
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Update/cr
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/$entry
      -- CP-element group 52: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/$entry
      -- 
    else_choice_transition_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_706_branch_ack_0, ack => sendB_CP_1657_elements(52)); -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(52), ack => type_cast_584_inst_req_0); -- 
    cr_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(52), ack => type_cast_584_inst_req_1); -- 
    -- CP-element group 53:  transition  output  delay-element  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	4 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	57 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 53: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/$exit
      -- CP-element group 53: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_582_konst_delay_trans
      -- CP-element group 53: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_req
      -- CP-element group 53: 	 branch_block_stmt_527/bbx_xnph_forx_xbody_PhiReq/phi_stmt_578/$exit
      -- 
    phi_stmt_578_req_2088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_578_req_2088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(53), ack => phi_stmt_578_req_0); -- 
    -- Element group sendB_CP_1657_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => sendB_CP_1657_elements(4), ack => sendB_CP_1657_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Sample/ra
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_0, ack => sendB_CP_1657_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	52 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (2) 
      -- CP-element group 55: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/Update/ca
      -- 
    ca_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_584_inst_ack_1, ack => sendB_CP_1657_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (6) 
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/$exit
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/$exit
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/$exit
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_sources/type_cast_584/SplitProtocol/$exit
      -- CP-element group 56: 	 branch_block_stmt_527/forx_xbody_forx_xbody_PhiReq/phi_stmt_578/phi_stmt_578_req
      -- 
    phi_stmt_578_req_2114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_578_req_2114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(56), ack => phi_stmt_578_req_1); -- 
    sendB_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "sendB_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendB_CP_1657_elements(54) & sendB_CP_1657_elements(55);
      gj_sendB_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendB_CP_1657_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  transition  place  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	53 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (2) 
      -- CP-element group 57: 	 branch_block_stmt_527/merge_stmt_577_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_527/merge_stmt_577_PhiAck/$entry
      -- 
    sendB_CP_1657_elements(57) <= OrReduce(sendB_CP_1657_elements(56) & sendB_CP_1657_elements(53));
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	5 
    -- CP-element group 58: 	6 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	18 
    -- CP-element group 58: 	20 
    -- CP-element group 58: 	22 
    -- CP-element group 58: 	24 
    -- CP-element group 58: 	8 
    -- CP-element group 58: 	12 
    -- CP-element group 58: 	26 
    -- CP-element group 58: 	10 
    -- CP-element group 58: 	14 
    -- CP-element group 58:  members (53) 
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/word_0/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_update_start
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/word_0/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_scale_1/scale_rename_req
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/merge_stmt_577__exit__
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_scale_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/word_access_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_scale_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Sample/req
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_scale_1/scale_rename_ack
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_resize_1/$exit
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_609_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_final_index_sum_regn_Update/req
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/ptr_deref_595_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_resize_1/index_resize_ack
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_complete/req
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_resize_1/index_resize_req
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_629_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_complete/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/addr_of_591_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_resize_1/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_619_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_computed_1
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_649_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_scaled_1
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705__entry__
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_599_update_start_
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/array_obj_ref_590_index_resized_1
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_659_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_639_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_527/assign_stmt_592_to_assign_stmt_705/type_cast_669_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_527/merge_stmt_577_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_527/merge_stmt_577_PhiAck/phi_stmt_578_ack
      -- 
    phi_stmt_578_ack_2119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_578_ack_0, ack => sendB_CP_1657_elements(58)); -- 
    cr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_609_inst_req_1); -- 
    cr_1835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_599_inst_req_1); -- 
    cr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1816_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => ptr_deref_595_load_0_req_1); -- 
    cr_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_649_inst_req_1); -- 
    req_1751_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1751_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => array_obj_ref_590_index_offset_req_0); -- 
    req_1756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => array_obj_ref_590_index_offset_req_1); -- 
    cr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_629_inst_req_1); -- 
    cr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_619_inst_req_1); -- 
    req_1771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => addr_of_591_final_reg_req_1); -- 
    cr_1891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_639_inst_req_1); -- 
    cr_1919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_659_inst_req_1); -- 
    cr_1933_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1933_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendB_CP_1657_elements(58), ack => type_cast_669_inst_req_1); -- 
    -- CP-element group 59:  merge  transition  place  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	2 
    -- CP-element group 59: 	51 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (16) 
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_716__exit__
      -- CP-element group 59: 	 branch_block_stmt_527/return__
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_714__exit__
      -- CP-element group 59: 	 branch_block_stmt_527/branch_block_stmt_527__exit__
      -- CP-element group 59: 	 branch_block_stmt_527/$exit
      -- CP-element group 59: 	 $exit
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_714_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_714_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_714_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_714_PhiAck/dummy
      -- CP-element group 59: 	 branch_block_stmt_527/return___PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_527/return___PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_716_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_716_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_716_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_527/merge_stmt_716_PhiAck/dummy
      -- 
    sendB_CP_1657_elements(59) <= OrReduce(sendB_CP_1657_elements(2) & sendB_CP_1657_elements(51));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_589_resized : std_logic_vector(13 downto 0);
    signal R_indvar_589_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_590_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_592 : std_logic_vector(31 downto 0);
    signal cmp68_533 : std_logic_vector(0 downto 0);
    signal conv12_610 : std_logic_vector(7 downto 0);
    signal conv18_620 : std_logic_vector(7 downto 0);
    signal conv24_630 : std_logic_vector(7 downto 0);
    signal conv30_640 : std_logic_vector(7 downto 0);
    signal conv36_650 : std_logic_vector(7 downto 0);
    signal conv42_660 : std_logic_vector(7 downto 0);
    signal conv48_670 : std_logic_vector(7 downto 0);
    signal conv_600 : std_logic_vector(7 downto 0);
    signal exitcond1_705 : std_logic_vector(0 downto 0);
    signal iNsTr_1_562 : std_logic_vector(63 downto 0);
    signal indvar_578 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_700 : std_logic_vector(63 downto 0);
    signal ptr_deref_595_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_595_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_595_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_595_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_595_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr15_616 : std_logic_vector(63 downto 0);
    signal shr21_626 : std_logic_vector(63 downto 0);
    signal shr27_636 : std_logic_vector(63 downto 0);
    signal shr33_646 : std_logic_vector(63 downto 0);
    signal shr39_656 : std_logic_vector(63 downto 0);
    signal shr45_666 : std_logic_vector(63 downto 0);
    signal shr9_606 : std_logic_vector(63 downto 0);
    signal shr_546 : std_logic_vector(31 downto 0);
    signal shrx_xop_558 : std_logic_vector(31 downto 0);
    signal tmp4_596 : std_logic_vector(63 downto 0);
    signal tmp72_575 : std_logic_vector(63 downto 0);
    signal tmp_552 : std_logic_vector(0 downto 0);
    signal type_cast_531_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_544_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_550_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_556_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_566_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_573_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_582_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_584_wire : std_logic_vector(63 downto 0);
    signal type_cast_604_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_614_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_634_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_644_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_654_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_698_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_568 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_590_constant_part_of_offset <= "00000000000000";
    array_obj_ref_590_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_590_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_590_resized_base_address <= "00000000000000";
    ptr_deref_595_word_offset_0 <= "00000000000000";
    type_cast_531_wire_constant <= "00000000000000000000000000000111";
    type_cast_544_wire_constant <= "00000000000000000000000000000011";
    type_cast_550_wire_constant <= "00000000000000000000000000000001";
    type_cast_556_wire_constant <= "11111111111111111111111111111111";
    type_cast_566_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_573_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_582_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_604_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_614_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_634_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_644_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_654_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_664_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_578: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_582_wire_constant & type_cast_584_wire;
      req <= phi_stmt_578_req_0 & phi_stmt_578_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_578",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_578_ack_0,
          idata => idata,
          odata => indvar_578,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_578
    -- flow-through select operator MUX_574_inst
    tmp72_575 <= xx_xop_568 when (tmp_552(0) /=  '0') else type_cast_573_wire_constant;
    addr_of_591_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_591_final_reg_req_0;
      addr_of_591_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_591_final_reg_req_1;
      addr_of_591_final_reg_ack_1<= rack(0);
      addr_of_591_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_591_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_590_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_592,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_561_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_561_inst_req_0;
      type_cast_561_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_561_inst_req_1;
      type_cast_561_inst_ack_1<= rack(0);
      type_cast_561_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_561_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shrx_xop_558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_1_562,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_584_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_584_inst_req_0;
      type_cast_584_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_584_inst_req_1;
      type_cast_584_inst_ack_1<= rack(0);
      type_cast_584_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_584_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_700,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_584_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_599_inst_req_0;
      type_cast_599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_599_inst_req_1;
      type_cast_599_inst_ack_1<= rack(0);
      type_cast_599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp4_596,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_609_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_609_inst_req_0;
      type_cast_609_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_609_inst_req_1;
      type_cast_609_inst_ack_1<= rack(0);
      type_cast_609_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_609_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr9_606,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_610,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_619_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_619_inst_req_0;
      type_cast_619_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_619_inst_req_1;
      type_cast_619_inst_ack_1<= rack(0);
      type_cast_619_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_619_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr15_616,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_620,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_629_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_629_inst_req_0;
      type_cast_629_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_629_inst_req_1;
      type_cast_629_inst_ack_1<= rack(0);
      type_cast_629_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_629_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr21_626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_639_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_639_inst_req_0;
      type_cast_639_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_639_inst_req_1;
      type_cast_639_inst_ack_1<= rack(0);
      type_cast_639_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_639_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr27_636,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_640,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_649_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_649_inst_req_0;
      type_cast_649_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_649_inst_req_1;
      type_cast_649_inst_ack_1<= rack(0);
      type_cast_649_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_649_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr33_646,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv36_650,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_659_inst_req_0;
      type_cast_659_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_659_inst_req_1;
      type_cast_659_inst_ack_1<= rack(0);
      type_cast_659_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_659_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr39_656,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv42_660,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_669_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_669_inst_req_0;
      type_cast_669_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_669_inst_req_1;
      type_cast_669_inst_ack_1<= rack(0);
      type_cast_669_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_669_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr45_666,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv48_670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_590_index_1_rename
    process(R_indvar_589_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_589_resized;
      ov(13 downto 0) := iv;
      R_indvar_589_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_590_index_1_resize
    process(indvar_578) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_578;
      ov := iv(13 downto 0);
      R_indvar_589_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_590_root_address_inst
    process(array_obj_ref_590_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_590_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_590_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_addr_0
    process(ptr_deref_595_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_595_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_595_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_base_resize
    process(arrayidx_592) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_592;
      ov := iv(13 downto 0);
      ptr_deref_595_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_gather_scatter
    process(ptr_deref_595_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_595_data_0;
      ov(63 downto 0) := iv;
      tmp4_596 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_595_root_address_inst
    process(ptr_deref_595_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_595_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_595_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_534_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp68_533;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_534_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_534_branch_req_0,
          ack0 => if_stmt_534_branch_ack_0,
          ack1 => if_stmt_534_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_706_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_705;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_706_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_706_branch_req_0,
          ack0 => if_stmt_706_branch_ack_0,
          ack1 => if_stmt_706_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_557_inst
    process(shr_546) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(shr_546, type_cast_556_wire_constant, tmp_var);
      shrx_xop_558 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_567_inst
    process(iNsTr_1_562) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_1_562, type_cast_566_wire_constant, tmp_var);
      xx_xop_568 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_699_inst
    process(indvar_578) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_578, type_cast_698_wire_constant, tmp_var);
      indvarx_xnext_700 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_704_inst
    process(indvarx_xnext_700, tmp72_575) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_700, tmp72_575, tmp_var);
      exitcond1_705 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_545_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(size_buffer, type_cast_544_wire_constant, tmp_var);
      shr_546 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_605_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_604_wire_constant, tmp_var);
      shr9_606 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_615_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_614_wire_constant, tmp_var);
      shr15_616 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_625_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_624_wire_constant, tmp_var);
      shr21_626 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_635_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_634_wire_constant, tmp_var);
      shr27_636 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_645_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_644_wire_constant, tmp_var);
      shr33_646 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_655_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_654_wire_constant, tmp_var);
      shr39_656 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_665_inst
    process(tmp4_596) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_596, type_cast_664_wire_constant, tmp_var);
      shr45_666 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_532_inst
    process(size_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(size_buffer, type_cast_531_wire_constant, tmp_var);
      cmp68_533 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_551_inst
    process(shr_546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(shr_546, type_cast_550_wire_constant, tmp_var);
      tmp_552 <= tmp_var; --
    end process;
    -- shared split operator group (14) : array_obj_ref_590_index_offset 
    ApIntAdd_group_14: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_589_scaled;
      array_obj_ref_590_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_590_index_offset_req_0;
      array_obj_ref_590_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_590_index_offset_req_1;
      array_obj_ref_590_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_14_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared load operator group (0) : ptr_deref_595_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_595_load_0_req_0;
      ptr_deref_595_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_595_load_0_req_1;
      ptr_deref_595_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_595_word_address_0;
      ptr_deref_595_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared outport operator group (0) : WPIPE_maxpool_output_pipe_671_inst WPIPE_maxpool_output_pipe_674_inst WPIPE_maxpool_output_pipe_677_inst WPIPE_maxpool_output_pipe_680_inst WPIPE_maxpool_output_pipe_683_inst WPIPE_maxpool_output_pipe_686_inst WPIPE_maxpool_output_pipe_689_inst WPIPE_maxpool_output_pipe_692_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_maxpool_output_pipe_671_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_maxpool_output_pipe_674_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_maxpool_output_pipe_677_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_maxpool_output_pipe_680_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_maxpool_output_pipe_683_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_maxpool_output_pipe_686_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_maxpool_output_pipe_689_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_maxpool_output_pipe_692_inst_req_0;
      WPIPE_maxpool_output_pipe_671_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_674_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_677_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_680_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_683_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_686_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_689_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_692_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_maxpool_output_pipe_671_inst_req_1;
      update_req_unguarded(6) <= WPIPE_maxpool_output_pipe_674_inst_req_1;
      update_req_unguarded(5) <= WPIPE_maxpool_output_pipe_677_inst_req_1;
      update_req_unguarded(4) <= WPIPE_maxpool_output_pipe_680_inst_req_1;
      update_req_unguarded(3) <= WPIPE_maxpool_output_pipe_683_inst_req_1;
      update_req_unguarded(2) <= WPIPE_maxpool_output_pipe_686_inst_req_1;
      update_req_unguarded(1) <= WPIPE_maxpool_output_pipe_689_inst_req_1;
      update_req_unguarded(0) <= WPIPE_maxpool_output_pipe_692_inst_req_1;
      WPIPE_maxpool_output_pipe_671_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_maxpool_output_pipe_674_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_maxpool_output_pipe_677_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_maxpool_output_pipe_680_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_maxpool_output_pipe_683_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_maxpool_output_pipe_686_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_maxpool_output_pipe_689_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_maxpool_output_pipe_692_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv48_670 & conv42_660 & conv36_650 & conv30_640 & conv24_630 & conv18_620 & conv12_610 & conv_600;
      maxpool_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "maxpool_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      maxpool_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "maxpool_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => maxpool_output_pipe_pipe_write_req(0),
          oack => maxpool_output_pipe_pipe_write_ack(0),
          odata => maxpool_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendModule is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
    output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
    output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendModule;
architecture sendModule_arch of sendModule is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendModule_CP_6819_start: Boolean;
  signal sendModule_CP_6819_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_3365_index_offset_req_0 : boolean;
  signal array_obj_ref_3365_index_offset_ack_1 : boolean;
  signal SUB_u16_u16_3278_inst_req_0 : boolean;
  signal n_row_3305_3268_buf_ack_0 : boolean;
  signal phi_stmt_3264_req_1 : boolean;
  signal phi_stmt_3259_ack_0 : boolean;
  signal SUB_u16_u16_3278_inst_ack_0 : boolean;
  signal type_cast_3252_inst_req_1 : boolean;
  signal n_row_3305_3268_buf_req_1 : boolean;
  signal type_cast_3252_inst_ack_0 : boolean;
  signal array_obj_ref_3365_index_offset_ack_0 : boolean;
  signal type_cast_3252_inst_req_0 : boolean;
  signal type_cast_3252_inst_ack_1 : boolean;
  signal n_col_3294_3263_buf_ack_1 : boolean;
  signal phi_stmt_3254_req_1 : boolean;
  signal phi_stmt_3264_req_0 : boolean;
  signal phi_stmt_3254_req_0 : boolean;
  signal phi_stmt_3254_ack_0 : boolean;
  signal ptr_deref_3380_load_0_ack_1 : boolean;
  signal n_row_3305_3268_buf_ack_1 : boolean;
  signal addr_of_3366_final_reg_req_0 : boolean;
  signal type_cast_3325_inst_req_0 : boolean;
  signal W_output_data1_3431_delayed_13_0_3558_inst_ack_0 : boolean;
  signal ptr_deref_3380_load_0_req_0 : boolean;
  signal W_output_data2_3455_delayed_13_0_3600_inst_ack_0 : boolean;
  signal SUB_u16_u16_3278_inst_req_1 : boolean;
  signal EQ_u3_u1_3668_inst_ack_1 : boolean;
  signal W_output_data2_3495_delayed_13_0_3670_inst_ack_0 : boolean;
  signal addr_of_3376_final_reg_req_1 : boolean;
  signal W_output_data2_3479_delayed_13_0_3642_inst_req_0 : boolean;
  signal phi_stmt_3264_ack_0 : boolean;
  signal array_obj_ref_3375_index_offset_ack_1 : boolean;
  signal addr_of_3366_final_reg_ack_0 : boolean;
  signal type_cast_3316_inst_req_0 : boolean;
  signal type_cast_3316_inst_ack_1 : boolean;
  signal W_output_data1_3431_delayed_13_0_3558_inst_req_0 : boolean;
  signal SUB_u16_u16_3278_inst_ack_1 : boolean;
  signal ptr_deref_3380_load_0_ack_0 : boolean;
  signal array_obj_ref_3375_index_offset_req_0 : boolean;
  signal W_output_data2_3479_delayed_13_0_3642_inst_ack_0 : boolean;
  signal type_cast_3316_inst_ack_0 : boolean;
  signal array_obj_ref_3375_index_offset_ack_0 : boolean;
  signal addr_of_3376_final_reg_req_0 : boolean;
  signal n_chl_3313_3258_buf_req_0 : boolean;
  signal n_chl_3313_3258_buf_ack_0 : boolean;
  signal array_obj_ref_3365_index_offset_req_1 : boolean;
  signal EQ_u3_u1_3682_inst_req_1 : boolean;
  signal W_output_data2_3455_delayed_13_0_3600_inst_req_0 : boolean;
  signal n_chl_3313_3258_buf_req_1 : boolean;
  signal n_chl_3313_3258_buf_ack_1 : boolean;
  signal n_address2_3357_3253_buf_req_0 : boolean;
  signal ptr_deref_3380_load_0_req_1 : boolean;
  signal addr_of_3376_final_reg_ack_0 : boolean;
  signal n_address2_3357_3253_buf_ack_0 : boolean;
  signal addr_of_3376_final_reg_ack_1 : boolean;
  signal array_obj_ref_3375_index_offset_req_1 : boolean;
  signal n_address2_3357_3253_buf_ack_1 : boolean;
  signal n_col_3294_3263_buf_req_1 : boolean;
  signal phi_stmt_3259_req_0 : boolean;
  signal RPIPE_output_pipe_3228_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3228_inst_ack_0 : boolean;
  signal n_row_3305_3268_buf_req_0 : boolean;
  signal RPIPE_output_pipe_3228_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3228_inst_ack_1 : boolean;
  signal n_col_3294_3263_buf_ack_0 : boolean;
  signal n_col_3294_3263_buf_req_0 : boolean;
  signal RPIPE_output_pipe_3231_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3231_inst_ack_0 : boolean;
  signal n_address2_3357_3253_buf_req_1 : boolean;
  signal RPIPE_output_pipe_3231_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3231_inst_ack_1 : boolean;
  signal phi_stmt_3259_req_1 : boolean;
  signal type_cast_3325_inst_ack_1 : boolean;
  signal addr_of_3366_final_reg_ack_1 : boolean;
  signal RPIPE_output_pipe_3234_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3234_inst_ack_0 : boolean;
  signal addr_of_3366_final_reg_req_1 : boolean;
  signal RPIPE_output_pipe_3234_inst_req_1 : boolean;
  signal RPIPE_output_pipe_3234_inst_ack_1 : boolean;
  signal type_cast_3325_inst_req_1 : boolean;
  signal type_cast_3325_inst_ack_0 : boolean;
  signal W_output_data2_3455_delayed_13_0_3600_inst_req_1 : boolean;
  signal do_while_stmt_3242_branch_req_0 : boolean;
  signal W_output_data2_3479_delayed_13_0_3642_inst_req_1 : boolean;
  signal W_output_data2_3455_delayed_13_0_3600_inst_ack_1 : boolean;
  signal phi_stmt_3244_req_1 : boolean;
  signal W_output_data2_3503_delayed_13_0_3684_inst_req_0 : boolean;
  signal phi_stmt_3244_req_0 : boolean;
  signal EQ_u3_u1_3682_inst_ack_0 : boolean;
  signal phi_stmt_3244_ack_0 : boolean;
  signal EQ_u3_u1_3584_inst_req_0 : boolean;
  signal EQ_u3_u1_3584_inst_ack_0 : boolean;
  signal type_cast_3316_inst_req_1 : boolean;
  signal W_output_data2_3479_delayed_13_0_3642_inst_ack_1 : boolean;
  signal n_address1_3343_3248_buf_req_0 : boolean;
  signal n_address1_3343_3248_buf_ack_0 : boolean;
  signal n_address1_3343_3248_buf_req_1 : boolean;
  signal n_address1_3343_3248_buf_ack_1 : boolean;
  signal phi_stmt_3249_req_1 : boolean;
  signal phi_stmt_3249_req_0 : boolean;
  signal phi_stmt_3249_ack_0 : boolean;
  signal EQ_u3_u1_3570_inst_ack_0 : boolean;
  signal EQ_u3_u1_3570_inst_req_0 : boolean;
  signal EQ_u3_u1_3626_inst_ack_1 : boolean;
  signal ptr_deref_3384_load_0_req_0 : boolean;
  signal ptr_deref_3384_load_0_ack_0 : boolean;
  signal EQ_u3_u1_3626_inst_req_1 : boolean;
  signal ptr_deref_3384_load_0_req_1 : boolean;
  signal ptr_deref_3384_load_0_ack_1 : boolean;
  signal W_output_data1_3431_delayed_13_0_3558_inst_ack_1 : boolean;
  signal W_output_data2_3503_delayed_13_0_3684_inst_req_1 : boolean;
  signal EQ_u3_u1_3654_inst_ack_1 : boolean;
  signal RPIPE_output_pipe_3387_inst_req_0 : boolean;
  signal RPIPE_output_pipe_3387_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3387_inst_req_1 : boolean;
  signal EQ_u3_u1_3626_inst_ack_0 : boolean;
  signal RPIPE_output_pipe_3387_inst_ack_1 : boolean;
  signal W_output_data2_3495_delayed_13_0_3670_inst_req_0 : boolean;
  signal EQ_u3_u1_3682_inst_req_0 : boolean;
  signal EQ_u3_u1_3654_inst_req_1 : boolean;
  signal EQ_u3_u1_3668_inst_req_1 : boolean;
  signal slice_3391_inst_req_0 : boolean;
  signal EQ_u3_u1_3626_inst_req_0 : boolean;
  signal slice_3391_inst_ack_0 : boolean;
  signal slice_3391_inst_req_1 : boolean;
  signal slice_3391_inst_ack_1 : boolean;
  signal W_output_data2_3503_delayed_13_0_3684_inst_ack_0 : boolean;
  signal W_output_data2_3503_delayed_13_0_3684_inst_ack_1 : boolean;
  signal EQ_u3_u1_3598_inst_ack_1 : boolean;
  signal EQ_u3_u1_3640_inst_ack_1 : boolean;
  signal EQ_u3_u1_3598_inst_req_1 : boolean;
  signal EQ_u3_u1_3640_inst_req_1 : boolean;
  signal slice_3395_inst_req_0 : boolean;
  signal slice_3395_inst_ack_0 : boolean;
  signal EQ_u3_u1_3668_inst_ack_0 : boolean;
  signal slice_3395_inst_req_1 : boolean;
  signal slice_3395_inst_ack_1 : boolean;
  signal W_output_data2_3495_delayed_13_0_3670_inst_ack_1 : boolean;
  signal W_output_data2_3495_delayed_13_0_3670_inst_req_1 : boolean;
  signal EQ_u3_u1_3598_inst_ack_0 : boolean;
  signal EQ_u3_u1_3668_inst_req_0 : boolean;
  signal slice_3399_inst_req_0 : boolean;
  signal slice_3399_inst_ack_0 : boolean;
  signal slice_3399_inst_req_1 : boolean;
  signal slice_3399_inst_ack_1 : boolean;
  signal EQ_u3_u1_3640_inst_ack_0 : boolean;
  signal EQ_u3_u1_3654_inst_ack_0 : boolean;
  signal EQ_u3_u1_3598_inst_req_0 : boolean;
  signal slice_3403_inst_req_0 : boolean;
  signal W_output_data2_3463_delayed_13_0_3614_inst_ack_1 : boolean;
  signal slice_3403_inst_ack_0 : boolean;
  signal slice_3403_inst_req_1 : boolean;
  signal W_output_data2_3463_delayed_13_0_3614_inst_req_1 : boolean;
  signal slice_3403_inst_ack_1 : boolean;
  signal W_output_data1_3439_delayed_13_0_3572_inst_ack_1 : boolean;
  signal EQ_u3_u1_3640_inst_req_0 : boolean;
  signal W_output_data1_3439_delayed_13_0_3572_inst_req_1 : boolean;
  signal EQ_u3_u1_3654_inst_req_0 : boolean;
  signal EQ_u3_u1_3556_inst_ack_1 : boolean;
  signal slice_3407_inst_req_0 : boolean;
  signal slice_3407_inst_ack_0 : boolean;
  signal slice_3407_inst_req_1 : boolean;
  signal slice_3407_inst_ack_1 : boolean;
  signal W_output_data1_3439_delayed_13_0_3572_inst_ack_0 : boolean;
  signal EQ_u3_u1_3556_inst_req_1 : boolean;
  signal W_output_data2_3447_delayed_13_0_3586_inst_ack_1 : boolean;
  signal W_output_data2_3447_delayed_13_0_3586_inst_req_1 : boolean;
  signal W_output_data2_3463_delayed_13_0_3614_inst_ack_0 : boolean;
  signal slice_3411_inst_req_0 : boolean;
  signal W_output_data2_3463_delayed_13_0_3614_inst_req_0 : boolean;
  signal slice_3411_inst_ack_0 : boolean;
  signal slice_3411_inst_req_1 : boolean;
  signal slice_3411_inst_ack_1 : boolean;
  signal W_output_data1_3439_delayed_13_0_3572_inst_req_0 : boolean;
  signal EQ_u3_u1_3682_inst_ack_1 : boolean;
  signal W_output_data2_3447_delayed_13_0_3586_inst_ack_0 : boolean;
  signal W_output_data2_3487_delayed_13_0_3656_inst_ack_1 : boolean;
  signal slice_3415_inst_req_0 : boolean;
  signal slice_3415_inst_ack_0 : boolean;
  signal EQ_u3_u1_3556_inst_ack_0 : boolean;
  signal W_output_data2_3487_delayed_13_0_3656_inst_req_1 : boolean;
  signal slice_3415_inst_req_1 : boolean;
  signal slice_3415_inst_ack_1 : boolean;
  signal EQ_u3_u1_3556_inst_req_0 : boolean;
  signal W_output_data2_3471_delayed_13_0_3628_inst_ack_1 : boolean;
  signal W_output_data2_3447_delayed_13_0_3586_inst_req_0 : boolean;
  signal slice_3419_inst_req_0 : boolean;
  signal slice_3419_inst_ack_0 : boolean;
  signal slice_3419_inst_req_1 : boolean;
  signal EQ_u3_u1_3612_inst_ack_1 : boolean;
  signal slice_3419_inst_ack_1 : boolean;
  signal W_output_data2_3471_delayed_13_0_3628_inst_req_1 : boolean;
  signal EQ_u3_u1_3612_inst_req_1 : boolean;
  signal W_output_data2_3487_delayed_13_0_3656_inst_ack_0 : boolean;
  signal slice_3423_inst_req_0 : boolean;
  signal slice_3423_inst_ack_0 : boolean;
  signal W_output_data2_3487_delayed_13_0_3656_inst_req_0 : boolean;
  signal slice_3423_inst_req_1 : boolean;
  signal slice_3423_inst_ack_1 : boolean;
  signal EQ_u3_u1_3570_inst_ack_1 : boolean;
  signal W_output_data2_3471_delayed_13_0_3628_inst_ack_0 : boolean;
  signal EQ_u3_u1_3584_inst_ack_1 : boolean;
  signal EQ_u3_u1_3584_inst_req_1 : boolean;
  signal EQ_u3_u1_3612_inst_ack_0 : boolean;
  signal slice_3427_inst_req_0 : boolean;
  signal EQ_u3_u1_3612_inst_req_0 : boolean;
  signal slice_3427_inst_ack_0 : boolean;
  signal slice_3427_inst_req_1 : boolean;
  signal slice_3427_inst_ack_1 : boolean;
  signal EQ_u3_u1_3570_inst_req_1 : boolean;
  signal W_output_data2_3471_delayed_13_0_3628_inst_req_0 : boolean;
  signal W_output_data1_3431_delayed_13_0_3558_inst_req_1 : boolean;
  signal slice_3431_inst_req_0 : boolean;
  signal slice_3431_inst_ack_0 : boolean;
  signal slice_3431_inst_req_1 : boolean;
  signal slice_3431_inst_ack_1 : boolean;
  signal slice_3435_inst_req_0 : boolean;
  signal slice_3435_inst_ack_0 : boolean;
  signal slice_3435_inst_req_1 : boolean;
  signal slice_3435_inst_ack_1 : boolean;
  signal slice_3439_inst_req_0 : boolean;
  signal slice_3439_inst_ack_0 : boolean;
  signal slice_3439_inst_req_1 : boolean;
  signal slice_3439_inst_ack_1 : boolean;
  signal slice_3443_inst_req_0 : boolean;
  signal slice_3443_inst_ack_0 : boolean;
  signal slice_3443_inst_req_1 : boolean;
  signal slice_3443_inst_ack_1 : boolean;
  signal slice_3447_inst_req_0 : boolean;
  signal slice_3447_inst_ack_0 : boolean;
  signal slice_3447_inst_req_1 : boolean;
  signal slice_3447_inst_ack_1 : boolean;
  signal slice_3451_inst_req_0 : boolean;
  signal slice_3451_inst_ack_0 : boolean;
  signal slice_3451_inst_req_1 : boolean;
  signal slice_3451_inst_ack_1 : boolean;
  signal slice_3455_inst_req_0 : boolean;
  signal slice_3455_inst_ack_0 : boolean;
  signal slice_3455_inst_req_1 : boolean;
  signal slice_3455_inst_ack_1 : boolean;
  signal slice_3459_inst_req_0 : boolean;
  signal slice_3459_inst_ack_0 : boolean;
  signal slice_3459_inst_req_1 : boolean;
  signal slice_3459_inst_ack_1 : boolean;
  signal EQ_u3_u1_3472_inst_req_0 : boolean;
  signal EQ_u3_u1_3472_inst_ack_0 : boolean;
  signal EQ_u3_u1_3472_inst_req_1 : boolean;
  signal EQ_u3_u1_3472_inst_ack_1 : boolean;
  signal W_output_data1_3383_delayed_13_0_3474_inst_req_0 : boolean;
  signal W_output_data1_3383_delayed_13_0_3474_inst_ack_0 : boolean;
  signal W_output_data1_3383_delayed_13_0_3474_inst_req_1 : boolean;
  signal W_output_data1_3383_delayed_13_0_3474_inst_ack_1 : boolean;
  signal EQ_u3_u1_3486_inst_req_0 : boolean;
  signal EQ_u3_u1_3486_inst_ack_0 : boolean;
  signal EQ_u3_u1_3486_inst_req_1 : boolean;
  signal EQ_u3_u1_3486_inst_ack_1 : boolean;
  signal W_output_data1_3391_delayed_13_0_3488_inst_req_0 : boolean;
  signal W_output_data1_3391_delayed_13_0_3488_inst_ack_0 : boolean;
  signal W_output_data1_3391_delayed_13_0_3488_inst_req_1 : boolean;
  signal W_output_data1_3391_delayed_13_0_3488_inst_ack_1 : boolean;
  signal EQ_u3_u1_3500_inst_req_0 : boolean;
  signal EQ_u3_u1_3500_inst_ack_0 : boolean;
  signal EQ_u3_u1_3500_inst_req_1 : boolean;
  signal EQ_u3_u1_3500_inst_ack_1 : boolean;
  signal W_output_data1_3399_delayed_13_0_3502_inst_req_0 : boolean;
  signal W_output_data1_3399_delayed_13_0_3502_inst_ack_0 : boolean;
  signal W_output_data1_3399_delayed_13_0_3502_inst_req_1 : boolean;
  signal W_output_data1_3399_delayed_13_0_3502_inst_ack_1 : boolean;
  signal EQ_u3_u1_3514_inst_req_0 : boolean;
  signal EQ_u3_u1_3514_inst_ack_0 : boolean;
  signal EQ_u3_u1_3514_inst_req_1 : boolean;
  signal EQ_u3_u1_3514_inst_ack_1 : boolean;
  signal W_output_data1_3407_delayed_13_0_3516_inst_req_0 : boolean;
  signal W_output_data1_3407_delayed_13_0_3516_inst_ack_0 : boolean;
  signal W_output_data1_3407_delayed_13_0_3516_inst_req_1 : boolean;
  signal W_output_data1_3407_delayed_13_0_3516_inst_ack_1 : boolean;
  signal EQ_u3_u1_3528_inst_req_0 : boolean;
  signal EQ_u3_u1_3528_inst_ack_0 : boolean;
  signal EQ_u3_u1_3528_inst_req_1 : boolean;
  signal EQ_u3_u1_3528_inst_ack_1 : boolean;
  signal W_output_data1_3415_delayed_13_0_3530_inst_req_0 : boolean;
  signal W_output_data1_3415_delayed_13_0_3530_inst_ack_0 : boolean;
  signal W_output_data1_3415_delayed_13_0_3530_inst_req_1 : boolean;
  signal W_output_data1_3415_delayed_13_0_3530_inst_ack_1 : boolean;
  signal EQ_u3_u1_3542_inst_req_0 : boolean;
  signal EQ_u3_u1_3542_inst_ack_0 : boolean;
  signal EQ_u3_u1_3542_inst_req_1 : boolean;
  signal EQ_u3_u1_3542_inst_ack_1 : boolean;
  signal W_output_data1_3423_delayed_13_0_3544_inst_req_0 : boolean;
  signal W_output_data1_3423_delayed_13_0_3544_inst_ack_0 : boolean;
  signal W_output_data1_3423_delayed_13_0_3544_inst_req_1 : boolean;
  signal W_output_data1_3423_delayed_13_0_3544_inst_ack_1 : boolean;
  signal W_fetch_addr1_3507_delayed_8_0_3693_inst_req_0 : boolean;
  signal W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_0 : boolean;
  signal W_fetch_addr1_3507_delayed_8_0_3693_inst_req_1 : boolean;
  signal W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3712_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3712_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3712_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3712_inst_ack_1 : boolean;
  signal ptr_deref_3697_store_0_req_0 : boolean;
  signal ptr_deref_3697_store_0_ack_0 : boolean;
  signal ptr_deref_3697_store_0_req_1 : boolean;
  signal ptr_deref_3697_store_0_ack_1 : boolean;
  signal W_fetch_addr2_3525_delayed_8_0_3714_inst_req_0 : boolean;
  signal W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_0 : boolean;
  signal W_fetch_addr2_3525_delayed_8_0_3714_inst_req_1 : boolean;
  signal W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_1 : boolean;
  signal CONCAT_u32_u64_3733_inst_req_0 : boolean;
  signal CONCAT_u32_u64_3733_inst_ack_0 : boolean;
  signal CONCAT_u32_u64_3733_inst_req_1 : boolean;
  signal CONCAT_u32_u64_3733_inst_ack_1 : boolean;
  signal ptr_deref_3718_store_0_req_0 : boolean;
  signal ptr_deref_3718_store_0_ack_0 : boolean;
  signal ptr_deref_3718_store_0_req_1 : boolean;
  signal ptr_deref_3718_store_0_ack_1 : boolean;
  signal SUB_u16_u16_3738_inst_req_0 : boolean;
  signal SUB_u16_u16_3738_inst_ack_0 : boolean;
  signal SUB_u16_u16_3738_inst_req_1 : boolean;
  signal SUB_u16_u16_3738_inst_ack_1 : boolean;
  signal do_while_stmt_3242_branch_ack_0 : boolean;
  signal do_while_stmt_3242_branch_ack_1 : boolean;
  signal WPIPE_input_done_pipe_3750_inst_req_0 : boolean;
  signal WPIPE_input_done_pipe_3750_inst_ack_0 : boolean;
  signal WPIPE_input_done_pipe_3750_inst_req_1 : boolean;
  signal WPIPE_input_done_pipe_3750_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendModule_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendModule_CP_6819_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendModule_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_6819_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendModule_CP_6819_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendModule_CP_6819_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendModule_CP_6819: Block -- control-path 
    signal sendModule_CP_6819_elements: BooleanArray(391 downto 0);
    -- 
  begin -- 
    sendModule_CP_6819_elements(0) <= sendModule_CP_6819_start;
    sendModule_CP_6819_symbol <= sendModule_CP_6819_elements(391);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3226/$entry
      -- CP-element group 0: 	 branch_block_stmt_3226/branch_block_stmt_3226__entry__
      -- CP-element group 0: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241__entry__
      -- CP-element group 0: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/$entry
      -- CP-element group 0: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Sample/rr
      -- 
    rr_6843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(0), ack => RPIPE_output_pipe_3228_inst_req_0); -- 
    -- CP-element group 1:  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	389 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	390 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_3226/do_while_stmt_3242__exit__
      -- CP-element group 1: 	 branch_block_stmt_3226/assign_stmt_3752__entry__
      -- CP-element group 1: 	 branch_block_stmt_3226/assign_stmt_3752/$entry
      -- CP-element group 1: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Sample/req
      -- 
    req_8270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(1), ack => WPIPE_input_done_pipe_3750_inst_req_0); -- 
    sendModule_CP_6819_elements(1) <= sendModule_CP_6819_elements(389);
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_update_start_
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Sample/ra
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Update/cr
      -- 
    ra_6844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3228_inst_ack_0, ack => sendModule_CP_6819_elements(2)); -- 
    cr_6848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(2), ack => RPIPE_output_pipe_3228_inst_req_1); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3228_Update/ca
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Sample/rr
      -- 
    ca_6849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3228_inst_ack_1, ack => sendModule_CP_6819_elements(3)); -- 
    rr_6857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(3), ack => RPIPE_output_pipe_3231_inst_req_0); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_update_start_
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Update/cr
      -- 
    ra_6858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3231_inst_ack_0, ack => sendModule_CP_6819_elements(4)); -- 
    cr_6862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(4), ack => RPIPE_output_pipe_3231_inst_req_1); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3231_Update/ca
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Sample/rr
      -- 
    ca_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3231_inst_ack_1, ack => sendModule_CP_6819_elements(5)); -- 
    rr_6871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(5), ack => RPIPE_output_pipe_3234_inst_req_0); -- 
    -- CP-element group 6:  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_update_start_
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Sample/ra
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Update/cr
      -- 
    ra_6872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3234_inst_ack_0, ack => sendModule_CP_6819_elements(6)); -- 
    cr_6876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(6), ack => RPIPE_output_pipe_3234_inst_req_1); -- 
    -- CP-element group 7:  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241__exit__
      -- CP-element group 7: 	 branch_block_stmt_3226/do_while_stmt_3242__entry__
      -- CP-element group 7: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/$exit
      -- CP-element group 7: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_3226/assign_stmt_3229_to_assign_stmt_3241/RPIPE_output_pipe_3234_Update/ca
      -- 
    ca_6877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3234_inst_ack_1, ack => sendModule_CP_6819_elements(7)); -- 
    -- CP-element group 8:  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (2) 
      -- CP-element group 8: 	 branch_block_stmt_3226/do_while_stmt_3242/$entry
      -- CP-element group 8: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242__entry__
      -- 
    sendModule_CP_6819_elements(8) <= sendModule_CP_6819_elements(7);
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	389 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242__exit__
      -- 
    -- Element group sendModule_CP_6819_elements(9) is bound as output of CP function.
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	13 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_back
      -- 
    -- Element group sendModule_CP_6819_elements(10) is bound as output of CP function.
    -- CP-element group 11:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	387 
    -- CP-element group 11: 	388 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_3226/do_while_stmt_3242/condition_done
      -- CP-element group 11: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_exit/$entry
      -- CP-element group 11: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_taken/$entry
      -- 
    sendModule_CP_6819_elements(11) <= sendModule_CP_6819_elements(16);
    -- CP-element group 12:  branch  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	386 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_body_done
      -- 
    sendModule_CP_6819_elements(12) <= sendModule_CP_6819_elements(386);
    -- CP-element group 13:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	10 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	44 
    -- CP-element group 13: 	65 
    -- CP-element group 13: 	84 
    -- CP-element group 13: 	103 
    -- CP-element group 13: 	27 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/back_edge_to_loop_body
      -- 
    sendModule_CP_6819_elements(13) <= sendModule_CP_6819_elements(10);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	8 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	46 
    -- CP-element group 14: 	67 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	105 
    -- CP-element group 14: 	29 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/first_time_through_loop_body
      -- 
    sendModule_CP_6819_elements(14) <= sendModule_CP_6819_elements(8);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	116 
    -- CP-element group 15: 	120 
    -- CP-element group 15: 	124 
    -- CP-element group 15: 	129 
    -- CP-element group 15: 	130 
    -- CP-element group 15: 	136 
    -- CP-element group 15: 	137 
    -- CP-element group 15: 	150 
    -- CP-element group 15: 	378 
    -- CP-element group 15: 	382 
    -- CP-element group 15: 	40 
    -- CP-element group 15: 	41 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	79 
    -- CP-element group 15: 	97 
    -- CP-element group 15: 	98 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	22 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/$entry
      -- CP-element group 15: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/loop_body_start
      -- 
    -- Element group sendModule_CP_6819_elements(15) is bound as output of CP function.
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	119 
    -- CP-element group 16: 	381 
    -- CP-element group 16: 	382 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/condition_evaluated
      -- 
    condition_evaluated_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(16), ack => do_while_stmt_3242_branch_req_0); -- 
    sendModule_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 15);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(119) & sendModule_CP_6819_elements(381) & sendModule_CP_6819_elements(382) & sendModule_CP_6819_elements(20);
      gj_sendModule_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	40 
    -- CP-element group 17: 	59 
    -- CP-element group 17: 	78 
    -- CP-element group 17: 	97 
    -- CP-element group 17: 	21 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	61 
    -- CP-element group 17: 	80 
    -- CP-element group 17: 	99 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/aggregated_phi_sample_req
      -- CP-element group 17: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_sample_start__ps
      -- 
    sendModule_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(40) & sendModule_CP_6819_elements(59) & sendModule_CP_6819_elements(78) & sendModule_CP_6819_elements(97) & sendModule_CP_6819_elements(21) & sendModule_CP_6819_elements(20);
      gj_sendModule_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	42 
    -- CP-element group 18: 	62 
    -- CP-element group 18: 	81 
    -- CP-element group 18: 	100 
    -- CP-element group 18: 	24 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	117 
    -- CP-element group 18: 	121 
    -- CP-element group 18: 	125 
    -- CP-element group 18: 	386 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	40 
    -- CP-element group 18: 	59 
    -- CP-element group 18: 	78 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	21 
    -- CP-element group 18:  members (6) 
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/aggregated_phi_sample_ack
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_sample_completed_
      -- 
    sendModule_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(42) & sendModule_CP_6819_elements(62) & sendModule_CP_6819_elements(81) & sendModule_CP_6819_elements(100) & sendModule_CP_6819_elements(24);
      gj_sendModule_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	41 
    -- CP-element group 19: 	60 
    -- CP-element group 19: 	79 
    -- CP-element group 19: 	98 
    -- CP-element group 19: 	22 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	82 
    -- CP-element group 19: 	101 
    -- CP-element group 19: 	25 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/aggregated_phi_update_req
      -- CP-element group 19: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_update_start__ps
      -- 
    sendModule_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(41) & sendModule_CP_6819_elements(60) & sendModule_CP_6819_elements(79) & sendModule_CP_6819_elements(98) & sendModule_CP_6819_elements(22);
      gj_sendModule_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	43 
    -- CP-element group 20: 	64 
    -- CP-element group 20: 	83 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	26 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/aggregated_phi_update_ack
      -- 
    sendModule_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(64) & sendModule_CP_6819_elements(83) & sendModule_CP_6819_elements(102) & sendModule_CP_6819_elements(26);
      gj_sendModule_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	15 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	119 
    -- CP-element group 21: 	123 
    -- CP-element group 21: 	18 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_sample_start_
      -- 
    sendModule_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(119) & sendModule_CP_6819_elements(123) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	15 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	131 
    -- CP-element group 22: 	228 
    -- CP-element group 22: 	236 
    -- CP-element group 22: 	244 
    -- CP-element group 22: 	252 
    -- CP-element group 22: 	260 
    -- CP-element group 22: 	268 
    -- CP-element group 22: 	276 
    -- CP-element group 22: 	284 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	19 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_update_start_
      -- 
    sendModule_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(131) & sendModule_CP_6819_elements(228) & sendModule_CP_6819_elements(236) & sendModule_CP_6819_elements(244) & sendModule_CP_6819_elements(252) & sendModule_CP_6819_elements(260) & sendModule_CP_6819_elements(268) & sendModule_CP_6819_elements(276) & sendModule_CP_6819_elements(284);
      gj_sendModule_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_sample_start__ps
      -- 
    sendModule_CP_6819_elements(23) <= sendModule_CP_6819_elements(17);
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	18 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	19 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_update_start__ps
      -- 
    sendModule_CP_6819_elements(25) <= sendModule_CP_6819_elements(19);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	131 
    -- CP-element group 26: 	226 
    -- CP-element group 26: 	234 
    -- CP-element group 26: 	242 
    -- CP-element group 26: 	250 
    -- CP-element group 26: 	258 
    -- CP-element group 26: 	266 
    -- CP-element group 26: 	274 
    -- CP-element group 26: 	282 
    -- CP-element group 26: 	20 
    -- CP-element group 26:  members (15) 
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_computed_1
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_resize_1/$entry
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_resize_1/$exit
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_resize_1/index_resize_req
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_resize_1/index_resize_ack
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_scale_1/$entry
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_scale_1/scale_rename_req
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_scale_1/$exit
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_scale_1/scale_rename_ack
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_scaled_1
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_index_resized_1
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_update_completed__ps
      -- 
    req_7194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(26), ack => array_obj_ref_3365_index_offset_req_0); -- 
    -- Element group sendModule_CP_6819_elements(26) is bound as output of CP function.
    -- CP-element group 27:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	13 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_loopback_trigger
      -- 
    sendModule_CP_6819_elements(27) <= sendModule_CP_6819_elements(13);
    -- CP-element group 28:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_loopback_sample_req
      -- CP-element group 28: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_loopback_sample_req_ps
      -- 
    phi_stmt_3244_loopback_sample_req_6907_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3244_loopback_sample_req_6907_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(28), ack => phi_stmt_3244_req_1); -- 
    -- Element group sendModule_CP_6819_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	14 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_entry_trigger
      -- 
    sendModule_CP_6819_elements(29) <= sendModule_CP_6819_elements(14);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_entry_sample_req
      -- CP-element group 30: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_entry_sample_req_ps
      -- 
    phi_stmt_3244_entry_sample_req_6910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3244_entry_sample_req_6910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(30), ack => phi_stmt_3244_req_0); -- 
    -- Element group sendModule_CP_6819_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_phi_mux_ack
      -- CP-element group 31: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3244_phi_mux_ack_ps
      -- 
    phi_stmt_3244_phi_mux_ack_6913_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3244_ack_0, ack => sendModule_CP_6819_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_sample_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_update_start_
      -- 
    -- Element group sendModule_CP_6819_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_update_completed__ps
      -- 
    sendModule_CP_6819_elements(34) <= sendModule_CP_6819_elements(35);
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3247_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(33), ack => sendModule_CP_6819_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_sample_start__ps
      -- CP-element group 36: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Sample/req
      -- 
    req_6934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(36), ack => n_address1_3343_3248_buf_req_0); -- 
    -- Element group sendModule_CP_6819_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_update_start__ps
      -- CP-element group 37: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_update_start_
      -- CP-element group 37: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Update/req
      -- 
    req_6939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(37), ack => n_address1_3343_3248_buf_req_1); -- 
    -- Element group sendModule_CP_6819_elements(37) is bound as output of CP function.
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_sample_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Sample/ack
      -- 
    ack_6935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3343_3248_buf_ack_0, ack => sendModule_CP_6819_elements(38)); -- 
    -- CP-element group 39:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address1_3248_Update/ack
      -- 
    ack_6940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address1_3343_3248_buf_ack_1, ack => sendModule_CP_6819_elements(39)); -- 
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	15 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	119 
    -- CP-element group 40: 	127 
    -- CP-element group 40: 	18 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	17 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_sample_start_
      -- 
    sendModule_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(119) & sendModule_CP_6819_elements(127) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	15 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	138 
    -- CP-element group 41: 	292 
    -- CP-element group 41: 	300 
    -- CP-element group 41: 	308 
    -- CP-element group 41: 	316 
    -- CP-element group 41: 	324 
    -- CP-element group 41: 	332 
    -- CP-element group 41: 	340 
    -- CP-element group 41: 	348 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	19 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_update_start_
      -- 
    sendModule_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 1,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(138) & sendModule_CP_6819_elements(292) & sendModule_CP_6819_elements(300) & sendModule_CP_6819_elements(308) & sendModule_CP_6819_elements(316) & sendModule_CP_6819_elements(324) & sendModule_CP_6819_elements(332) & sendModule_CP_6819_elements(340) & sendModule_CP_6819_elements(348);
      gj_sendModule_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	18 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	138 
    -- CP-element group 43: 	290 
    -- CP-element group 43: 	298 
    -- CP-element group 43: 	306 
    -- CP-element group 43: 	314 
    -- CP-element group 43: 	322 
    -- CP-element group 43: 	330 
    -- CP-element group 43: 	338 
    -- CP-element group 43: 	346 
    -- CP-element group 43: 	20 
    -- CP-element group 43:  members (15) 
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_resized_1
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_scaled_1
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_resize_1/index_resize_req
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_computed_1
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_resize_1/index_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Sample/$entry
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_scale_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_scale_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_scale_1/scale_rename_req
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_scale_1/scale_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Sample/req
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_resize_1/$entry
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_index_resize_1/$exit
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_update_completed__ps
      -- 
    req_7240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(43), ack => array_obj_ref_3375_index_offset_req_0); -- 
    -- Element group sendModule_CP_6819_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	13 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_loopback_trigger
      -- 
    sendModule_CP_6819_elements(44) <= sendModule_CP_6819_elements(13);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_loopback_sample_req
      -- CP-element group 45: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_loopback_sample_req_ps
      -- 
    phi_stmt_3249_loopback_sample_req_6951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3249_loopback_sample_req_6951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(45), ack => phi_stmt_3249_req_1); -- 
    -- Element group sendModule_CP_6819_elements(45) is bound as output of CP function.
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	14 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_entry_trigger
      -- 
    sendModule_CP_6819_elements(46) <= sendModule_CP_6819_elements(14);
    -- CP-element group 47:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_entry_sample_req
      -- CP-element group 47: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_entry_sample_req_ps
      -- 
    phi_stmt_3249_entry_sample_req_6954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3249_entry_sample_req_6954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(47), ack => phi_stmt_3249_req_0); -- 
    -- Element group sendModule_CP_6819_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_phi_mux_ack
      -- CP-element group 48: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3249_phi_mux_ack_ps
      -- 
    phi_stmt_3249_phi_mux_ack_6957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3249_ack_0, ack => sendModule_CP_6819_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_sample_start__ps
      -- 
    -- Element group sendModule_CP_6819_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_update_start__ps
      -- 
    -- Element group sendModule_CP_6819_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	53 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Sample/rr
      -- CP-element group 51: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_sample_start_
      -- 
    rr_6970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(51), ack => type_cast_3252_inst_req_0); -- 
    sendModule_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(49) & sendModule_CP_6819_elements(53);
      gj_sendModule_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_update_start_
      -- CP-element group 52: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Update/cr
      -- 
    cr_6975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(52), ack => type_cast_3252_inst_req_1); -- 
    sendModule_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(50) & sendModule_CP_6819_elements(54);
      gj_sendModule_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	51 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Sample/ra
      -- CP-element group 53: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_sample_completed__ps
      -- 
    ra_6971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3252_inst_ack_0, ack => sendModule_CP_6819_elements(53)); -- 
    -- CP-element group 54:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_Update/ca
      -- CP-element group 54: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3252_update_completed__ps
      -- 
    ca_6976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3252_inst_ack_1, ack => sendModule_CP_6819_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Sample/req
      -- 
    req_6988_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6988_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(55), ack => n_address2_3357_3253_buf_req_0); -- 
    -- Element group sendModule_CP_6819_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_update_start_
      -- CP-element group 56: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Update/req
      -- 
    req_6993_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6993_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(56), ack => n_address2_3357_3253_buf_req_1); -- 
    -- Element group sendModule_CP_6819_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_sample_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_sample_completed_
      -- CP-element group 57: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Sample/ack
      -- 
    ack_6989_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3357_3253_buf_ack_0, ack => sendModule_CP_6819_elements(57)); -- 
    -- CP-element group 58:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (4) 
      -- CP-element group 58: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_update_completed__ps
      -- CP-element group 58: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Update/$exit
      -- CP-element group 58: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_address2_3253_Update/ack
      -- 
    ack_6994_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_address2_3357_3253_buf_ack_1, ack => sendModule_CP_6819_elements(58)); -- 
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	119 
    -- CP-element group 59: 	18 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	17 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_sample_start_
      -- 
    sendModule_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(119) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	15 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	64 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	19 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_update_start_
      -- 
    sendModule_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(64);
      gj_sendModule_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	17 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_sample_start__ps
      -- 
    sendModule_CP_6819_elements(61) <= sendModule_CP_6819_elements(17);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	18 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(62) is bound as output of CP function.
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_update_start__ps
      -- 
    sendModule_CP_6819_elements(63) <= sendModule_CP_6819_elements(19);
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	60 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_update_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(64) is bound as output of CP function.
    -- CP-element group 65:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	13 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_loopback_trigger
      -- 
    sendModule_CP_6819_elements(65) <= sendModule_CP_6819_elements(13);
    -- CP-element group 66:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (2) 
      -- CP-element group 66: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_loopback_sample_req
      -- CP-element group 66: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_loopback_sample_req_ps
      -- 
    phi_stmt_3254_loopback_sample_req_7005_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3254_loopback_sample_req_7005_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(66), ack => phi_stmt_3254_req_1); -- 
    -- Element group sendModule_CP_6819_elements(66) is bound as output of CP function.
    -- CP-element group 67:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	14 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_entry_trigger
      -- 
    sendModule_CP_6819_elements(67) <= sendModule_CP_6819_elements(14);
    -- CP-element group 68:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_entry_sample_req_ps
      -- CP-element group 68: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_entry_sample_req
      -- 
    phi_stmt_3254_entry_sample_req_7008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3254_entry_sample_req_7008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(68), ack => phi_stmt_3254_req_0); -- 
    -- Element group sendModule_CP_6819_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (2) 
      -- CP-element group 69: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_phi_mux_ack
      -- CP-element group 69: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3254_phi_mux_ack_ps
      -- 
    phi_stmt_3254_phi_mux_ack_7011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3254_ack_0, ack => sendModule_CP_6819_elements(69)); -- 
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_sample_start__ps
      -- CP-element group 70: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_sample_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (2) 
      -- CP-element group 71: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_update_start__ps
      -- CP-element group 71: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_update_start_
      -- 
    -- Element group sendModule_CP_6819_elements(71) is bound as output of CP function.
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	73 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_update_completed__ps
      -- 
    sendModule_CP_6819_elements(72) <= sendModule_CP_6819_elements(73);
    -- CP-element group 73:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	72 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3257_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(71), ack => sendModule_CP_6819_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_sample_start__ps
      -- CP-element group 74: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Sample/req
      -- 
    req_7032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(74), ack => n_chl_3313_3258_buf_req_0); -- 
    -- Element group sendModule_CP_6819_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_update_start__ps
      -- CP-element group 75: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_update_start_
      -- CP-element group 75: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Update/req
      -- 
    req_7037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(75), ack => n_chl_3313_3258_buf_req_1); -- 
    -- Element group sendModule_CP_6819_elements(75) is bound as output of CP function.
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_sample_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Sample/ack
      -- 
    ack_7033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3313_3258_buf_ack_0, ack => sendModule_CP_6819_elements(76)); -- 
    -- CP-element group 77:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (4) 
      -- CP-element group 77: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_chl_3258_Update/ack
      -- 
    ack_7038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_chl_3313_3258_buf_ack_1, ack => sendModule_CP_6819_elements(77)); -- 
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	18 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	17 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_sample_start_
      -- 
    sendModule_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	15 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	83 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	19 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_update_start_
      -- 
    sendModule_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(83);
      gj_sendModule_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	17 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_sample_start__ps
      -- 
    sendModule_CP_6819_elements(80) <= sendModule_CP_6819_elements(17);
    -- CP-element group 81:  join  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	18 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(81) is bound as output of CP function.
    -- CP-element group 82:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	19 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_update_start__ps
      -- 
    sendModule_CP_6819_elements(82) <= sendModule_CP_6819_elements(19);
    -- CP-element group 83:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	20 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	79 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_update_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(83) is bound as output of CP function.
    -- CP-element group 84:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	13 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_loopback_trigger
      -- 
    sendModule_CP_6819_elements(84) <= sendModule_CP_6819_elements(13);
    -- CP-element group 85:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_loopback_sample_req_ps
      -- CP-element group 85: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_loopback_sample_req
      -- 
    phi_stmt_3259_loopback_sample_req_7049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3259_loopback_sample_req_7049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(85), ack => phi_stmt_3259_req_1); -- 
    -- Element group sendModule_CP_6819_elements(85) is bound as output of CP function.
    -- CP-element group 86:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_entry_trigger
      -- 
    sendModule_CP_6819_elements(86) <= sendModule_CP_6819_elements(14);
    -- CP-element group 87:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_entry_sample_req_ps
      -- CP-element group 87: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_entry_sample_req
      -- 
    phi_stmt_3259_entry_sample_req_7052_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3259_entry_sample_req_7052_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(87), ack => phi_stmt_3259_req_0); -- 
    -- Element group sendModule_CP_6819_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_phi_mux_ack
      -- CP-element group 88: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3259_phi_mux_ack_ps
      -- 
    phi_stmt_3259_phi_mux_ack_7055_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3259_ack_0, ack => sendModule_CP_6819_elements(88)); -- 
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_sample_start_
      -- CP-element group 89: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_sample_start__ps
      -- CP-element group 89: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_update_start_
      -- CP-element group 90: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_update_start__ps
      -- 
    -- Element group sendModule_CP_6819_elements(90) is bound as output of CP function.
    -- CP-element group 91:  join  transition  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: successors 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_update_completed__ps
      -- 
    sendModule_CP_6819_elements(91) <= sendModule_CP_6819_elements(92);
    -- CP-element group 92:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (1) 
      -- CP-element group 92: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3262_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(90), ack => sendModule_CP_6819_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_sample_start__ps
      -- CP-element group 93: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_sample_start_
      -- CP-element group 93: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Sample/req
      -- CP-element group 93: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Sample/$entry
      -- 
    req_7076_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7076_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(93), ack => n_col_3294_3263_buf_req_0); -- 
    -- Element group sendModule_CP_6819_elements(93) is bound as output of CP function.
    -- CP-element group 94:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	96 
    -- CP-element group 94:  members (4) 
      -- CP-element group 94: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_update_start_
      -- CP-element group 94: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_update_start__ps
      -- CP-element group 94: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Update/req
      -- CP-element group 94: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Update/$entry
      -- 
    req_7081_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7081_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(94), ack => n_col_3294_3263_buf_req_1); -- 
    -- Element group sendModule_CP_6819_elements(94) is bound as output of CP function.
    -- CP-element group 95:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (4) 
      -- CP-element group 95: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_sample_completed__ps
      -- CP-element group 95: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Sample/ack
      -- CP-element group 95: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Sample/$exit
      -- 
    ack_7077_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3294_3263_buf_ack_0, ack => sendModule_CP_6819_elements(95)); -- 
    -- CP-element group 96:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	94 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (4) 
      -- CP-element group 96: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Update/ack
      -- CP-element group 96: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_update_completed__ps
      -- CP-element group 96: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_col_3263_update_completed_
      -- 
    ack_7082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_col_3294_3263_buf_ack_1, ack => sendModule_CP_6819_elements(96)); -- 
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	15 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	119 
    -- CP-element group 97: 	18 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	17 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_sample_start_
      -- 
    sendModule_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(119) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  join  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	15 
    -- CP-element group 98: marked-predecessors 
    -- CP-element group 98: 	102 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	19 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_update_start_
      -- 
    sendModule_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendModule_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(102);
      gj_sendModule_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	17 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (1) 
      -- CP-element group 99: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_sample_start__ps
      -- 
    sendModule_CP_6819_elements(99) <= sendModule_CP_6819_elements(17);
    -- CP-element group 100:  join  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	18 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_sample_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(100) is bound as output of CP function.
    -- CP-element group 101:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	19 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_update_start__ps
      -- 
    sendModule_CP_6819_elements(101) <= sendModule_CP_6819_elements(19);
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: marked-successors 
    -- CP-element group 102: 	98 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_update_completed__ps
      -- 
    -- Element group sendModule_CP_6819_elements(102) is bound as output of CP function.
    -- CP-element group 103:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	13 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (1) 
      -- CP-element group 103: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_loopback_trigger
      -- 
    sendModule_CP_6819_elements(103) <= sendModule_CP_6819_elements(13);
    -- CP-element group 104:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_loopback_sample_req
      -- CP-element group 104: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_loopback_sample_req_ps
      -- 
    phi_stmt_3264_loopback_sample_req_7093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3264_loopback_sample_req_7093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(104), ack => phi_stmt_3264_req_1); -- 
    -- Element group sendModule_CP_6819_elements(104) is bound as output of CP function.
    -- CP-element group 105:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	14 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_entry_trigger
      -- 
    sendModule_CP_6819_elements(105) <= sendModule_CP_6819_elements(14);
    -- CP-element group 106:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_entry_sample_req_ps
      -- CP-element group 106: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_entry_sample_req
      -- 
    phi_stmt_3264_entry_sample_req_7096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3264_entry_sample_req_7096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(106), ack => phi_stmt_3264_req_0); -- 
    -- Element group sendModule_CP_6819_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_phi_mux_ack
      -- CP-element group 107: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/phi_stmt_3264_phi_mux_ack_ps
      -- 
    phi_stmt_3264_phi_mux_ack_7099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3264_ack_0, ack => sendModule_CP_6819_elements(107)); -- 
    -- CP-element group 108:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (4) 
      -- CP-element group 108: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_sample_start__ps
      -- CP-element group 108: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_sample_completed__ps
      -- CP-element group 108: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_sample_start_
      -- 
    -- Element group sendModule_CP_6819_elements(108) is bound as output of CP function.
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_update_start__ps
      -- CP-element group 109: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_update_start_
      -- 
    -- Element group sendModule_CP_6819_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	111 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_update_completed__ps
      -- 
    sendModule_CP_6819_elements(110) <= sendModule_CP_6819_elements(111);
    -- CP-element group 111:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	110 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3267_update_completed_
      -- 
    -- Element group sendModule_CP_6819_elements(111) is a control-delay.
    cp_element_111_delay: control_delay_element  generic map(name => " 111_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(109), ack => sendModule_CP_6819_elements(111), clk => clk, reset =>reset);
    -- CP-element group 112:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (4) 
      -- CP-element group 112: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Sample/req
      -- CP-element group 112: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_sample_start__ps
      -- 
    req_7120_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7120_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(112), ack => n_row_3305_3268_buf_req_0); -- 
    -- Element group sendModule_CP_6819_elements(112) is bound as output of CP function.
    -- CP-element group 113:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (4) 
      -- CP-element group 113: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_update_start_
      -- CP-element group 113: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Update/req
      -- CP-element group 113: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Update/$entry
      -- CP-element group 113: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_update_start__ps
      -- 
    req_7125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(113), ack => n_row_3305_3268_buf_req_1); -- 
    -- Element group sendModule_CP_6819_elements(113) is bound as output of CP function.
    -- CP-element group 114:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114:  members (4) 
      -- CP-element group 114: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_sample_completed__ps
      -- 
    ack_7121_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3305_3268_buf_ack_0, ack => sendModule_CP_6819_elements(114)); -- 
    -- CP-element group 115:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (4) 
      -- CP-element group 115: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_update_completed__ps
      -- CP-element group 115: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_Update/ack
      -- CP-element group 115: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/R_n_row_3268_update_completed_
      -- 
    ack_7126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_row_3305_3268_buf_ack_1, ack => sendModule_CP_6819_elements(115)); -- 
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	15 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	118 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Sample/$entry
      -- 
    rr_7135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(116), ack => SUB_u16_u16_3278_inst_req_0); -- 
    sendModule_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(118);
      gj_sendModule_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	18 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Update/$entry
      -- CP-element group 117: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Update/cr
      -- CP-element group 117: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_update_start_
      -- 
    cr_7140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(117), ack => SUB_u16_u16_3278_inst_req_1); -- 
    sendModule_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(18) & sendModule_CP_6819_elements(119);
      gj_sendModule_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: marked-successors 
    -- CP-element group 118: 	116 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Sample/$exit
      -- CP-element group 118: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Sample/ra
      -- CP-element group 118: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_sample_completed_
      -- 
    ra_7136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3278_inst_ack_0, ack => sendModule_CP_6819_elements(118)); -- 
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	16 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	40 
    -- CP-element group 119: 	59 
    -- CP-element group 119: 	97 
    -- CP-element group 119: 	21 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Update/$exit
      -- CP-element group 119: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_Update/ca
      -- CP-element group 119: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3278_update_completed_
      -- 
    ca_7141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3278_inst_ack_1, ack => sendModule_CP_6819_elements(119)); -- 
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	15 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	122 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Sample/rr
      -- CP-element group 120: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_sample_start_
      -- CP-element group 120: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Sample/$entry
      -- 
    rr_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(120), ack => type_cast_3316_inst_req_0); -- 
    sendModule_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(122);
      gj_sendModule_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	18 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_update_start_
      -- CP-element group 121: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Update/cr
      -- 
    cr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(121), ack => type_cast_3316_inst_req_1); -- 
    sendModule_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(18) & sendModule_CP_6819_elements(123);
      gj_sendModule_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: marked-successors 
    -- CP-element group 122: 	120 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Sample/$exit
      -- CP-element group 122: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Sample/ra
      -- CP-element group 122: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_sample_completed_
      -- 
    ra_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3316_inst_ack_0, ack => sendModule_CP_6819_elements(122)); -- 
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	386 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	21 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Update/$exit
      -- CP-element group 123: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_Update/ca
      -- CP-element group 123: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3316_update_completed_
      -- 
    ca_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3316_inst_ack_1, ack => sendModule_CP_6819_elements(123)); -- 
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	15 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	126 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Sample/rr
      -- CP-element group 124: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_sample_start_
      -- CP-element group 124: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Sample/$entry
      -- 
    rr_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(124), ack => type_cast_3325_inst_req_0); -- 
    sendModule_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(126);
      gj_sendModule_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	18 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_update_start_
      -- CP-element group 125: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Update/cr
      -- CP-element group 125: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Update/$entry
      -- 
    cr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(125), ack => type_cast_3325_inst_req_1); -- 
    sendModule_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(18) & sendModule_CP_6819_elements(127);
      gj_sendModule_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: marked-successors 
    -- CP-element group 126: 	124 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_sample_completed_
      -- CP-element group 126: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Sample/ra
      -- 
    ra_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3325_inst_ack_0, ack => sendModule_CP_6819_elements(126)); -- 
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	386 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: 	40 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_update_completed_
      -- CP-element group 127: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Update/ca
      -- CP-element group 127: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/type_cast_3325_Update/$exit
      -- 
    ca_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3325_inst_ack_1, ack => sendModule_CP_6819_elements(127)); -- 
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	132 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	133 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_request/$entry
      -- CP-element group 128: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_request/req
      -- CP-element group 128: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_sample_start_
      -- 
    req_7209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(128), ack => addr_of_3366_final_reg_req_0); -- 
    sendModule_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(132) & sendModule_CP_6819_elements(133);
      gj_sendModule_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	15 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	144 
    -- CP-element group 129: 	356 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	134 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_complete/$entry
      -- CP-element group 129: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_update_start_
      -- CP-element group 129: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_complete/req
      -- 
    req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(129), ack => addr_of_3366_final_reg_req_1); -- 
    sendModule_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(144) & sendModule_CP_6819_elements(356);
      gj_sendModule_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	15 
    -- CP-element group 130: marked-predecessors 
    -- CP-element group 130: 	133 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	132 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_update_start
      -- CP-element group 130: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Update/req
      -- 
    req_7199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(130), ack => array_obj_ref_3365_index_offset_req_1); -- 
    sendModule_cp_element_group_130: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_130"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(133);
      gj_sendModule_cp_element_group_130 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(130), clk => clk, reset => reset); --
    end block;
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	26 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	386 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	22 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Sample/ack
      -- CP-element group 131: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_sample_complete
      -- CP-element group 131: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Sample/$exit
      -- 
    ack_7195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3365_index_offset_ack_0, ack => sendModule_CP_6819_elements(131)); -- 
    -- CP-element group 132:  transition  input  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	130 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	128 
    -- CP-element group 132:  members (8) 
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Update/ack
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_base_plus_offset/sum_rename_ack
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_final_index_sum_regn_Update/$exit
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_base_plus_offset/$entry
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_base_plus_offset/$exit
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_base_plus_offset/sum_rename_req
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_offset_calculated
      -- CP-element group 132: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3365_root_address_calculated
      -- 
    ack_7200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3365_index_offset_ack_1, ack => sendModule_CP_6819_elements(132)); -- 
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	130 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_request/$exit
      -- CP-element group 133: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_request/ack
      -- CP-element group 133: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_sample_completed_
      -- 
    ack_7210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3366_final_reg_ack_0, ack => sendModule_CP_6819_elements(133)); -- 
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	129 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	142 
    -- CP-element group 134: 	354 
    -- CP-element group 134:  members (19) 
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_address_resized
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_word_addrgen/root_register_ack
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_addr_resize/$entry
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_addr_resize/$exit
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_addr_resize/base_resize_req
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_addr_resize/base_resize_ack
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_word_addrgen/root_register_req
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_plus_offset/$entry
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_plus_offset/$exit
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_plus_offset/sum_rename_req
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_base_plus_offset/sum_rename_ack
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_word_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_word_addrgen/$entry
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_word_addrgen/$exit
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_root_address_calculated
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_complete/$exit
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3366_complete/ack
      -- 
    ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3366_final_reg_ack_1, ack => sendModule_CP_6819_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	139 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	140 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	140 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_request/$entry
      -- CP-element group 135: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_request/req
      -- CP-element group 135: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_sample_start_
      -- 
    req_7255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(135), ack => addr_of_3376_final_reg_req_0); -- 
    sendModule_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(139) & sendModule_CP_6819_elements(140);
      gj_sendModule_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	15 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	148 
    -- CP-element group 136: 	368 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	141 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_complete/$entry
      -- CP-element group 136: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_complete/req
      -- CP-element group 136: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_update_start_
      -- 
    req_7260_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7260_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(136), ack => addr_of_3376_final_reg_req_1); -- 
    sendModule_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(148) & sendModule_CP_6819_elements(368);
      gj_sendModule_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	15 
    -- CP-element group 137: marked-predecessors 
    -- CP-element group 137: 	140 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	139 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_update_start
      -- CP-element group 137: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Update/req
      -- 
    req_7245_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7245_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(137), ack => array_obj_ref_3375_index_offset_req_1); -- 
    sendModule_cp_element_group_137: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_137"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(140);
      gj_sendModule_cp_element_group_137 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(137), clk => clk, reset => reset); --
    end block;
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	43 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	386 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	41 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Sample/ack
      -- CP-element group 138: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_sample_complete
      -- 
    ack_7241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3375_index_offset_ack_0, ack => sendModule_CP_6819_elements(138)); -- 
    -- CP-element group 139:  transition  input  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	137 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	135 
    -- CP-element group 139:  members (8) 
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_base_plus_offset/sum_rename_ack
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_base_plus_offset/$entry
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_base_plus_offset/$exit
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_root_address_calculated
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Update/ack
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_offset_calculated
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_final_index_sum_regn_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/array_obj_ref_3375_base_plus_offset/sum_rename_req
      -- 
    ack_7246_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3375_index_offset_ack_1, ack => sendModule_CP_6819_elements(139)); -- 
    -- CP-element group 140:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: successors 
    -- CP-element group 140: marked-successors 
    -- CP-element group 140: 	135 
    -- CP-element group 140: 	137 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_request/$exit
      -- CP-element group 140: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_request/ack
      -- CP-element group 140: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_sample_completed_
      -- 
    ack_7256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3376_final_reg_ack_0, ack => sendModule_CP_6819_elements(140)); -- 
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	136 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	146 
    -- CP-element group 141: 	366 
    -- CP-element group 141:  members (19) 
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_complete/$exit
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_word_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_root_address_calculated
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_complete/ack
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/addr_of_3376_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_address_resized
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_addr_resize/$entry
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_addr_resize/$exit
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_addr_resize/base_resize_req
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_addr_resize/base_resize_ack
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_plus_offset/$entry
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_plus_offset/$exit
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_plus_offset/sum_rename_req
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_base_plus_offset/sum_rename_ack
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_word_addrgen/$entry
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_word_addrgen/$exit
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_word_addrgen/root_register_req
      -- CP-element group 141: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_word_addrgen/root_register_ack
      -- 
    ack_7261_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3376_final_reg_ack_1, ack => sendModule_CP_6819_elements(141)); -- 
    -- CP-element group 142:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	134 
    -- CP-element group 142: marked-predecessors 
    -- CP-element group 142: 	376 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	144 
    -- CP-element group 142:  members (5) 
      -- CP-element group 142: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/$entry
      -- CP-element group 142: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_sample_start_
      -- CP-element group 142: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/word_0/rr
      -- CP-element group 142: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/$entry
      -- CP-element group 142: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/word_0/$entry
      -- 
    rr_7294_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7294_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(142), ack => ptr_deref_3380_load_0_req_0); -- 
    sendModule_cp_element_group_142: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_142"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(134) & sendModule_CP_6819_elements(376);
      gj_sendModule_cp_element_group_142 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(142), clk => clk, reset => reset); --
    end block;
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	164 
    -- CP-element group 143: 	168 
    -- CP-element group 143: 	172 
    -- CP-element group 143: 	176 
    -- CP-element group 143: 	180 
    -- CP-element group 143: 	184 
    -- CP-element group 143: 	188 
    -- CP-element group 143: 	192 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/$entry
      -- CP-element group 143: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/$entry
      -- CP-element group 143: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_update_start_
      -- CP-element group 143: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/word_0/cr
      -- 
    cr_7305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(143), ack => ptr_deref_3380_load_0_req_1); -- 
    sendModule_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(164) & sendModule_CP_6819_elements(168) & sendModule_CP_6819_elements(172) & sendModule_CP_6819_elements(176) & sendModule_CP_6819_elements(180) & sendModule_CP_6819_elements(184) & sendModule_CP_6819_elements(188) & sendModule_CP_6819_elements(192);
      gj_sendModule_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	142 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	383 
    -- CP-element group 144: marked-successors 
    -- CP-element group 144: 	129 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/$exit
      -- CP-element group 144: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/word_0/ra
      -- CP-element group 144: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Sample/word_access_start/word_0/$exit
      -- 
    ra_7295_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3380_load_0_ack_0, ack => sendModule_CP_6819_elements(144)); -- 
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145: 	166 
    -- CP-element group 145: 	170 
    -- CP-element group 145: 	174 
    -- CP-element group 145: 	178 
    -- CP-element group 145: 	182 
    -- CP-element group 145: 	186 
    -- CP-element group 145: 	190 
    -- CP-element group 145:  members (9) 
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/$exit
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/ptr_deref_3380_Merge/merge_ack
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/word_0/ca
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/ptr_deref_3380_Merge/$exit
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/ptr_deref_3380_Merge/merge_req
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/word_access_complete/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_Update/ptr_deref_3380_Merge/$entry
      -- 
    ca_7306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3380_load_0_ack_1, ack => sendModule_CP_6819_elements(145)); -- 
    -- CP-element group 146:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	141 
    -- CP-element group 146: marked-predecessors 
    -- CP-element group 146: 	376 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	148 
    -- CP-element group 146:  members (5) 
      -- CP-element group 146: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_sample_start_
      -- CP-element group 146: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/$entry
      -- CP-element group 146: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/$entry
      -- CP-element group 146: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/word_0/$entry
      -- CP-element group 146: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/word_0/rr
      -- 
    rr_7344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(146), ack => ptr_deref_3384_load_0_req_0); -- 
    sendModule_cp_element_group_146: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_146"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(141) & sendModule_CP_6819_elements(376);
      gj_sendModule_cp_element_group_146 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(146), clk => clk, reset => reset); --
    end block;
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	196 
    -- CP-element group 147: 	200 
    -- CP-element group 147: 	204 
    -- CP-element group 147: 	208 
    -- CP-element group 147: 	212 
    -- CP-element group 147: 	216 
    -- CP-element group 147: 	220 
    -- CP-element group 147: 	224 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (5) 
      -- CP-element group 147: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_update_start_
      -- CP-element group 147: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/$entry
      -- CP-element group 147: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/$entry
      -- CP-element group 147: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/word_0/$entry
      -- CP-element group 147: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/word_0/cr
      -- 
    cr_7355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(147), ack => ptr_deref_3384_load_0_req_1); -- 
    sendModule_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(196) & sendModule_CP_6819_elements(200) & sendModule_CP_6819_elements(204) & sendModule_CP_6819_elements(208) & sendModule_CP_6819_elements(212) & sendModule_CP_6819_elements(216) & sendModule_CP_6819_elements(220) & sendModule_CP_6819_elements(224);
      gj_sendModule_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	146 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	384 
    -- CP-element group 148: marked-successors 
    -- CP-element group 148: 	136 
    -- CP-element group 148:  members (5) 
      -- CP-element group 148: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/$exit
      -- CP-element group 148: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/word_0/$exit
      -- CP-element group 148: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Sample/word_access_start/word_0/ra
      -- 
    ra_7345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3384_load_0_ack_0, ack => sendModule_CP_6819_elements(148)); -- 
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	194 
    -- CP-element group 149: 	198 
    -- CP-element group 149: 	202 
    -- CP-element group 149: 	206 
    -- CP-element group 149: 	210 
    -- CP-element group 149: 	214 
    -- CP-element group 149: 	218 
    -- CP-element group 149: 	222 
    -- CP-element group 149:  members (9) 
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/$exit
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/word_0/$exit
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/word_access_complete/word_0/ca
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/ptr_deref_3384_Merge/$entry
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/ptr_deref_3384_Merge/$exit
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/ptr_deref_3384_Merge/merge_req
      -- CP-element group 149: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_Update/ptr_deref_3384_Merge/merge_ack
      -- 
    ca_7356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3384_load_0_ack_1, ack => sendModule_CP_6819_elements(149)); -- 
    -- CP-element group 150:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	15 
    -- CP-element group 150: marked-predecessors 
    -- CP-element group 150: 	153 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	152 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_sample_start_
      -- CP-element group 150: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Sample/$entry
      -- CP-element group 150: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Sample/rr
      -- 
    rr_7369_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7369_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(150), ack => RPIPE_output_pipe_3387_inst_req_0); -- 
    sendModule_cp_element_group_150: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_150"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(153);
      gj_sendModule_cp_element_group_150 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(150), clk => clk, reset => reset); --
    end block;
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	156 
    -- CP-element group 151: 	160 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_update_start_
      -- CP-element group 151: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Update/$entry
      -- CP-element group 151: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Update/cr
      -- 
    cr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(151), ack => RPIPE_output_pipe_3387_inst_req_1); -- 
    sendModule_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(152) & sendModule_CP_6819_elements(156) & sendModule_CP_6819_elements(160);
      gj_sendModule_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  transition  input  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	150 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	151 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Sample/ra
      -- 
    ra_7370_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3387_inst_ack_0, ack => sendModule_CP_6819_elements(152)); -- 
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	154 
    -- CP-element group 153: 	158 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	150 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/RPIPE_output_pipe_3387_Update/ca
      -- 
    ca_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_output_pipe_3387_inst_ack_1, ack => sendModule_CP_6819_elements(153)); -- 
    -- CP-element group 154:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	153 
    -- CP-element group 154: marked-predecessors 
    -- CP-element group 154: 	156 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	156 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_sample_start_
      -- CP-element group 154: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Sample/$entry
      -- CP-element group 154: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Sample/rr
      -- 
    rr_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(154), ack => slice_3391_inst_req_0); -- 
    sendModule_cp_element_group_154: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_154"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(153) & sendModule_CP_6819_elements(156);
      gj_sendModule_cp_element_group_154 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(154), clk => clk, reset => reset); --
    end block;
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	232 
    -- CP-element group 155: 	240 
    -- CP-element group 155: 	248 
    -- CP-element group 155: 	256 
    -- CP-element group 155: 	264 
    -- CP-element group 155: 	272 
    -- CP-element group 155: 	280 
    -- CP-element group 155: 	288 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_update_start_
      -- CP-element group 155: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Update/$entry
      -- CP-element group 155: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Update/cr
      -- 
    cr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(155), ack => slice_3391_inst_req_1); -- 
    sendModule_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(232) & sendModule_CP_6819_elements(240) & sendModule_CP_6819_elements(248) & sendModule_CP_6819_elements(256) & sendModule_CP_6819_elements(264) & sendModule_CP_6819_elements(272) & sendModule_CP_6819_elements(280) & sendModule_CP_6819_elements(288);
      gj_sendModule_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	154 
    -- CP-element group 156: successors 
    -- CP-element group 156: marked-successors 
    -- CP-element group 156: 	151 
    -- CP-element group 156: 	154 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Sample/ra
      -- 
    ra_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3391_inst_ack_0, ack => sendModule_CP_6819_elements(156)); -- 
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	230 
    -- CP-element group 157: 	238 
    -- CP-element group 157: 	246 
    -- CP-element group 157: 	254 
    -- CP-element group 157: 	262 
    -- CP-element group 157: 	270 
    -- CP-element group 157: 	278 
    -- CP-element group 157: 	286 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3391_Update/ca
      -- 
    ca_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3391_inst_ack_1, ack => sendModule_CP_6819_elements(157)); -- 
    -- CP-element group 158:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	153 
    -- CP-element group 158: marked-predecessors 
    -- CP-element group 158: 	160 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	160 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_sample_start_
      -- CP-element group 158: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Sample/$entry
      -- CP-element group 158: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Sample/rr
      -- 
    rr_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(158), ack => slice_3395_inst_req_0); -- 
    sendModule_cp_element_group_158: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_158"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(153) & sendModule_CP_6819_elements(160);
      gj_sendModule_cp_element_group_158 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(158), clk => clk, reset => reset); --
    end block;
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	296 
    -- CP-element group 159: 	304 
    -- CP-element group 159: 	312 
    -- CP-element group 159: 	320 
    -- CP-element group 159: 	328 
    -- CP-element group 159: 	336 
    -- CP-element group 159: 	344 
    -- CP-element group 159: 	352 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_update_start_
      -- CP-element group 159: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Update/$entry
      -- CP-element group 159: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Update/cr
      -- 
    cr_7402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(159), ack => slice_3395_inst_req_1); -- 
    sendModule_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(296) & sendModule_CP_6819_elements(304) & sendModule_CP_6819_elements(312) & sendModule_CP_6819_elements(320) & sendModule_CP_6819_elements(328) & sendModule_CP_6819_elements(336) & sendModule_CP_6819_elements(344) & sendModule_CP_6819_elements(352);
      gj_sendModule_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	158 
    -- CP-element group 160: successors 
    -- CP-element group 160: marked-successors 
    -- CP-element group 160: 	151 
    -- CP-element group 160: 	158 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Sample/ra
      -- 
    ra_7398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3395_inst_ack_0, ack => sendModule_CP_6819_elements(160)); -- 
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	294 
    -- CP-element group 161: 	302 
    -- CP-element group 161: 	310 
    -- CP-element group 161: 	318 
    -- CP-element group 161: 	326 
    -- CP-element group 161: 	334 
    -- CP-element group 161: 	342 
    -- CP-element group 161: 	350 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3395_Update/ca
      -- 
    ca_7403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3395_inst_ack_1, ack => sendModule_CP_6819_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	145 
    -- CP-element group 162: marked-predecessors 
    -- CP-element group 162: 	164 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	164 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Sample/rr
      -- 
    rr_7411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(162), ack => slice_3399_inst_req_0); -- 
    sendModule_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(164);
      gj_sendModule_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	360 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_update_start_
      -- CP-element group 163: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Update/$entry
      -- CP-element group 163: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Update/cr
      -- 
    cr_7416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(163), ack => slice_3399_inst_req_1); -- 
    sendModule_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	162 
    -- CP-element group 164: successors 
    -- CP-element group 164: marked-successors 
    -- CP-element group 164: 	143 
    -- CP-element group 164: 	162 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_sample_completed_
      -- CP-element group 164: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Sample/$exit
      -- CP-element group 164: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Sample/ra
      -- 
    ra_7412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3399_inst_ack_0, ack => sendModule_CP_6819_elements(164)); -- 
    -- CP-element group 165:  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	358 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_update_completed_
      -- CP-element group 165: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Update/$exit
      -- CP-element group 165: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3399_Update/ca
      -- 
    ca_7417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3399_inst_ack_1, ack => sendModule_CP_6819_elements(165)); -- 
    -- CP-element group 166:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	145 
    -- CP-element group 166: marked-predecessors 
    -- CP-element group 166: 	168 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	168 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_sample_start_
      -- CP-element group 166: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Sample/$entry
      -- CP-element group 166: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Sample/rr
      -- 
    rr_7425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(166), ack => slice_3403_inst_req_0); -- 
    sendModule_cp_element_group_166: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_166"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(168);
      gj_sendModule_cp_element_group_166 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(166), clk => clk, reset => reset); --
    end block;
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	360 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_update_start_
      -- CP-element group 167: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Update/cr
      -- 
    cr_7430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(167), ack => slice_3403_inst_req_1); -- 
    sendModule_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	166 
    -- CP-element group 168: successors 
    -- CP-element group 168: marked-successors 
    -- CP-element group 168: 	143 
    -- CP-element group 168: 	166 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Sample/ra
      -- 
    ra_7426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3403_inst_ack_0, ack => sendModule_CP_6819_elements(168)); -- 
    -- CP-element group 169:  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	358 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3403_Update/ca
      -- 
    ca_7431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3403_inst_ack_1, ack => sendModule_CP_6819_elements(169)); -- 
    -- CP-element group 170:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	145 
    -- CP-element group 170: marked-predecessors 
    -- CP-element group 170: 	172 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	172 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_sample_start_
      -- CP-element group 170: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Sample/$entry
      -- CP-element group 170: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Sample/rr
      -- 
    rr_7439_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7439_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(170), ack => slice_3407_inst_req_0); -- 
    sendModule_cp_element_group_170: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_170"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(172);
      gj_sendModule_cp_element_group_170 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(170), clk => clk, reset => reset); --
    end block;
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	360 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_update_start_
      -- CP-element group 171: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Update/$entry
      -- CP-element group 171: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Update/cr
      -- 
    cr_7444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(171), ack => slice_3407_inst_req_1); -- 
    sendModule_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	170 
    -- CP-element group 172: successors 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	143 
    -- CP-element group 172: 	170 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Sample/ra
      -- 
    ra_7440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3407_inst_ack_0, ack => sendModule_CP_6819_elements(172)); -- 
    -- CP-element group 173:  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	358 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3407_Update/ca
      -- 
    ca_7445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3407_inst_ack_1, ack => sendModule_CP_6819_elements(173)); -- 
    -- CP-element group 174:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	145 
    -- CP-element group 174: marked-predecessors 
    -- CP-element group 174: 	176 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	176 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_sample_start_
      -- CP-element group 174: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Sample/$entry
      -- CP-element group 174: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Sample/rr
      -- 
    rr_7453_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7453_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(174), ack => slice_3411_inst_req_0); -- 
    sendModule_cp_element_group_174: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_174"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(176);
      gj_sendModule_cp_element_group_174 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(174), clk => clk, reset => reset); --
    end block;
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	360 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_update_start_
      -- CP-element group 175: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Update/$entry
      -- CP-element group 175: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Update/cr
      -- 
    cr_7458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(175), ack => slice_3411_inst_req_1); -- 
    sendModule_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	174 
    -- CP-element group 176: successors 
    -- CP-element group 176: marked-successors 
    -- CP-element group 176: 	143 
    -- CP-element group 176: 	174 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Sample/ra
      -- 
    ra_7454_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3411_inst_ack_0, ack => sendModule_CP_6819_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	358 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3411_Update/ca
      -- 
    ca_7459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3411_inst_ack_1, ack => sendModule_CP_6819_elements(177)); -- 
    -- CP-element group 178:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	145 
    -- CP-element group 178: marked-predecessors 
    -- CP-element group 178: 	180 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	180 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_sample_start_
      -- CP-element group 178: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Sample/$entry
      -- CP-element group 178: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Sample/rr
      -- 
    rr_7467_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7467_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(178), ack => slice_3415_inst_req_0); -- 
    sendModule_cp_element_group_178: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_178"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(180);
      gj_sendModule_cp_element_group_178 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(178), clk => clk, reset => reset); --
    end block;
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	360 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_update_start_
      -- CP-element group 179: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Update/$entry
      -- CP-element group 179: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Update/cr
      -- 
    cr_7472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(179), ack => slice_3415_inst_req_1); -- 
    sendModule_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	178 
    -- CP-element group 180: successors 
    -- CP-element group 180: marked-successors 
    -- CP-element group 180: 	143 
    -- CP-element group 180: 	178 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Sample/ra
      -- 
    ra_7468_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3415_inst_ack_0, ack => sendModule_CP_6819_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	358 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3415_Update/ca
      -- 
    ca_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3415_inst_ack_1, ack => sendModule_CP_6819_elements(181)); -- 
    -- CP-element group 182:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	145 
    -- CP-element group 182: marked-predecessors 
    -- CP-element group 182: 	184 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	184 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_sample_start_
      -- CP-element group 182: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Sample/$entry
      -- CP-element group 182: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Sample/rr
      -- 
    rr_7481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(182), ack => slice_3419_inst_req_0); -- 
    sendModule_cp_element_group_182: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_182"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(184);
      gj_sendModule_cp_element_group_182 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(182), clk => clk, reset => reset); --
    end block;
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	360 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_update_start_
      -- CP-element group 183: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Update/$entry
      -- CP-element group 183: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Update/cr
      -- 
    cr_7486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(183), ack => slice_3419_inst_req_1); -- 
    sendModule_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	182 
    -- CP-element group 184: successors 
    -- CP-element group 184: marked-successors 
    -- CP-element group 184: 	143 
    -- CP-element group 184: 	182 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Sample/ra
      -- 
    ra_7482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3419_inst_ack_0, ack => sendModule_CP_6819_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	358 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3419_Update/ca
      -- 
    ca_7487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3419_inst_ack_1, ack => sendModule_CP_6819_elements(185)); -- 
    -- CP-element group 186:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	145 
    -- CP-element group 186: marked-predecessors 
    -- CP-element group 186: 	188 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	188 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_sample_start_
      -- CP-element group 186: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Sample/$entry
      -- CP-element group 186: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Sample/rr
      -- 
    rr_7495_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7495_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(186), ack => slice_3423_inst_req_0); -- 
    sendModule_cp_element_group_186: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_186"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(188);
      gj_sendModule_cp_element_group_186 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(186), clk => clk, reset => reset); --
    end block;
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	360 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_update_start_
      -- CP-element group 187: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Update/$entry
      -- CP-element group 187: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Update/cr
      -- 
    cr_7500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(187), ack => slice_3423_inst_req_1); -- 
    sendModule_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	186 
    -- CP-element group 188: successors 
    -- CP-element group 188: marked-successors 
    -- CP-element group 188: 	143 
    -- CP-element group 188: 	186 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Sample/ra
      -- 
    ra_7496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3423_inst_ack_0, ack => sendModule_CP_6819_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	358 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_update_completed_
      -- CP-element group 189: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3423_Update/ca
      -- 
    ca_7501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3423_inst_ack_1, ack => sendModule_CP_6819_elements(189)); -- 
    -- CP-element group 190:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	145 
    -- CP-element group 190: marked-predecessors 
    -- CP-element group 190: 	192 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	192 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_sample_start_
      -- CP-element group 190: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Sample/$entry
      -- CP-element group 190: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Sample/rr
      -- 
    rr_7509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(190), ack => slice_3427_inst_req_0); -- 
    sendModule_cp_element_group_190: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_190"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(145) & sendModule_CP_6819_elements(192);
      gj_sendModule_cp_element_group_190 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(190), clk => clk, reset => reset); --
    end block;
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	360 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_update_start_
      -- CP-element group 191: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Update/$entry
      -- CP-element group 191: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Update/cr
      -- 
    cr_7514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(191), ack => slice_3427_inst_req_1); -- 
    sendModule_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	190 
    -- CP-element group 192: successors 
    -- CP-element group 192: marked-successors 
    -- CP-element group 192: 	143 
    -- CP-element group 192: 	190 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Sample/ra
      -- 
    ra_7510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3427_inst_ack_0, ack => sendModule_CP_6819_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	358 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Update/$exit
      -- CP-element group 193: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3427_Update/ca
      -- 
    ca_7515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3427_inst_ack_1, ack => sendModule_CP_6819_elements(193)); -- 
    -- CP-element group 194:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	149 
    -- CP-element group 194: marked-predecessors 
    -- CP-element group 194: 	196 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	196 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_sample_start_
      -- CP-element group 194: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Sample/$entry
      -- CP-element group 194: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Sample/rr
      -- 
    rr_7523_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7523_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(194), ack => slice_3431_inst_req_0); -- 
    sendModule_cp_element_group_194: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_194"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(196);
      gj_sendModule_cp_element_group_194 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(194), clk => clk, reset => reset); --
    end block;
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	372 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	197 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_update_start_
      -- CP-element group 195: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Update/$entry
      -- CP-element group 195: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Update/cr
      -- 
    cr_7528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(195), ack => slice_3431_inst_req_1); -- 
    sendModule_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	194 
    -- CP-element group 196: successors 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	147 
    -- CP-element group 196: 	194 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Sample/ra
      -- 
    ra_7524_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3431_inst_ack_0, ack => sendModule_CP_6819_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	195 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	370 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3431_Update/ca
      -- 
    ca_7529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3431_inst_ack_1, ack => sendModule_CP_6819_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	149 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Sample/$entry
      -- CP-element group 198: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Sample/rr
      -- 
    rr_7537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(198), ack => slice_3435_inst_req_0); -- 
    sendModule_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(200);
      gj_sendModule_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	372 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_update_start_
      -- CP-element group 199: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Update/$entry
      -- CP-element group 199: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Update/cr
      -- 
    cr_7542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(199), ack => slice_3435_inst_req_1); -- 
    sendModule_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	147 
    -- CP-element group 200: 	198 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Sample/ra
      -- 
    ra_7538_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3435_inst_ack_0, ack => sendModule_CP_6819_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	370 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_update_completed_
      -- CP-element group 201: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3435_Update/ca
      -- 
    ca_7543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3435_inst_ack_1, ack => sendModule_CP_6819_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	149 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Sample/rr
      -- 
    rr_7551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(202), ack => slice_3439_inst_req_0); -- 
    sendModule_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(204);
      gj_sendModule_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	372 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_update_start_
      -- CP-element group 203: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Update/cr
      -- 
    cr_7556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(203), ack => slice_3439_inst_req_1); -- 
    sendModule_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	147 
    -- CP-element group 204: 	202 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Sample/ra
      -- 
    ra_7552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3439_inst_ack_0, ack => sendModule_CP_6819_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	370 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3439_Update/ca
      -- 
    ca_7557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3439_inst_ack_1, ack => sendModule_CP_6819_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	149 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Sample/rr
      -- 
    rr_7565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(206), ack => slice_3443_inst_req_0); -- 
    sendModule_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(208);
      gj_sendModule_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	372 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_update_start_
      -- CP-element group 207: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Update/cr
      -- 
    cr_7570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(207), ack => slice_3443_inst_req_1); -- 
    sendModule_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	147 
    -- CP-element group 208: 	206 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Sample/ra
      -- 
    ra_7566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3443_inst_ack_0, ack => sendModule_CP_6819_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	370 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3443_Update/ca
      -- 
    ca_7571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3443_inst_ack_1, ack => sendModule_CP_6819_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	149 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Sample/rr
      -- 
    rr_7579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(210), ack => slice_3447_inst_req_0); -- 
    sendModule_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(212);
      gj_sendModule_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	372 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_update_start_
      -- CP-element group 211: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Update/cr
      -- 
    cr_7584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(211), ack => slice_3447_inst_req_1); -- 
    sendModule_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	147 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Sample/ra
      -- 
    ra_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3447_inst_ack_0, ack => sendModule_CP_6819_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	370 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3447_Update/ca
      -- 
    ca_7585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3447_inst_ack_1, ack => sendModule_CP_6819_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	149 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Sample/rr
      -- 
    rr_7593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(214), ack => slice_3451_inst_req_0); -- 
    sendModule_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(216);
      gj_sendModule_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	372 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_update_start_
      -- CP-element group 215: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Update/cr
      -- 
    cr_7598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(215), ack => slice_3451_inst_req_1); -- 
    sendModule_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	147 
    -- CP-element group 216: 	214 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Sample/ra
      -- 
    ra_7594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3451_inst_ack_0, ack => sendModule_CP_6819_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	370 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3451_Update/ca
      -- 
    ca_7599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3451_inst_ack_1, ack => sendModule_CP_6819_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	149 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Sample/rr
      -- 
    rr_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(218), ack => slice_3455_inst_req_0); -- 
    sendModule_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(220);
      gj_sendModule_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	372 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_update_start_
      -- CP-element group 219: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Update/cr
      -- 
    cr_7612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(219), ack => slice_3455_inst_req_1); -- 
    sendModule_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	147 
    -- CP-element group 220: 	218 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Sample/ra
      -- 
    ra_7608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3455_inst_ack_0, ack => sendModule_CP_6819_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	370 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3455_Update/ca
      -- 
    ca_7613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3455_inst_ack_1, ack => sendModule_CP_6819_elements(221)); -- 
    -- CP-element group 222:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	149 
    -- CP-element group 222: marked-predecessors 
    -- CP-element group 222: 	224 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	224 
    -- CP-element group 222:  members (3) 
      -- CP-element group 222: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_sample_start_
      -- CP-element group 222: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Sample/$entry
      -- CP-element group 222: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Sample/rr
      -- 
    rr_7621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(222), ack => slice_3459_inst_req_0); -- 
    sendModule_cp_element_group_222: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_222"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(149) & sendModule_CP_6819_elements(224);
      gj_sendModule_cp_element_group_222 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(222), clk => clk, reset => reset); --
    end block;
    -- CP-element group 223:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: marked-predecessors 
    -- CP-element group 223: 	372 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	225 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_update_start_
      -- CP-element group 223: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Update/$entry
      -- CP-element group 223: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Update/cr
      -- 
    cr_7626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(223), ack => slice_3459_inst_req_1); -- 
    sendModule_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	222 
    -- CP-element group 224: successors 
    -- CP-element group 224: marked-successors 
    -- CP-element group 224: 	147 
    -- CP-element group 224: 	222 
    -- CP-element group 224:  members (3) 
      -- CP-element group 224: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_sample_completed_
      -- CP-element group 224: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Sample/$exit
      -- CP-element group 224: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Sample/ra
      -- 
    ra_7622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3459_inst_ack_0, ack => sendModule_CP_6819_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	223 
    -- CP-element group 225: successors 
    -- CP-element group 225: 	370 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_update_completed_
      -- CP-element group 225: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Update/$exit
      -- CP-element group 225: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/slice_3459_Update/ca
      -- 
    ca_7627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_3459_inst_ack_1, ack => sendModule_CP_6819_elements(225)); -- 
    -- CP-element group 226:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	26 
    -- CP-element group 226: marked-predecessors 
    -- CP-element group 226: 	228 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	228 
    -- CP-element group 226:  members (3) 
      -- CP-element group 226: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Sample/rr
      -- 
    rr_7635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(226), ack => EQ_u3_u1_3472_inst_req_0); -- 
    sendModule_cp_element_group_226: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_226"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(228);
      gj_sendModule_cp_element_group_226 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(226), clk => clk, reset => reset); --
    end block;
    -- CP-element group 227:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: marked-predecessors 
    -- CP-element group 227: 	360 
    -- CP-element group 227: successors 
    -- CP-element group 227: 	229 
    -- CP-element group 227:  members (3) 
      -- CP-element group 227: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_update_start_
      -- CP-element group 227: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Update/$entry
      -- CP-element group 227: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Update/cr
      -- 
    cr_7640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(227), ack => EQ_u3_u1_3472_inst_req_1); -- 
    sendModule_cp_element_group_227: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_227"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_227 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(227), clk => clk, reset => reset); --
    end block;
    -- CP-element group 228:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: successors 
    -- CP-element group 228: marked-successors 
    -- CP-element group 228: 	226 
    -- CP-element group 228: 	22 
    -- CP-element group 228:  members (3) 
      -- CP-element group 228: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_sample_completed_
      -- CP-element group 228: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Sample/$exit
      -- CP-element group 228: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Sample/ra
      -- 
    ra_7636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3472_inst_ack_0, ack => sendModule_CP_6819_elements(228)); -- 
    -- CP-element group 229:  transition  input  bypass  pipeline-parent 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	227 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	358 
    -- CP-element group 229:  members (3) 
      -- CP-element group 229: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_update_completed_
      -- CP-element group 229: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Update/$exit
      -- CP-element group 229: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3472_Update/ca
      -- 
    ca_7641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 229_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3472_inst_ack_1, ack => sendModule_CP_6819_elements(229)); -- 
    -- CP-element group 230:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	157 
    -- CP-element group 230: marked-predecessors 
    -- CP-element group 230: 	232 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	232 
    -- CP-element group 230:  members (3) 
      -- CP-element group 230: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_sample_start_
      -- CP-element group 230: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Sample/$entry
      -- CP-element group 230: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Sample/req
      -- 
    req_7649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(230), ack => W_output_data1_3383_delayed_13_0_3474_inst_req_0); -- 
    sendModule_cp_element_group_230: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_230"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(232);
      gj_sendModule_cp_element_group_230 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(230), clk => clk, reset => reset); --
    end block;
    -- CP-element group 231:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: marked-predecessors 
    -- CP-element group 231: 	360 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	233 
    -- CP-element group 231:  members (3) 
      -- CP-element group 231: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_update_start_
      -- CP-element group 231: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Update/req
      -- 
    req_7654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(231), ack => W_output_data1_3383_delayed_13_0_3474_inst_req_1); -- 
    sendModule_cp_element_group_231: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_231"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_231 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(231), clk => clk, reset => reset); --
    end block;
    -- CP-element group 232:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	230 
    -- CP-element group 232: successors 
    -- CP-element group 232: marked-successors 
    -- CP-element group 232: 	155 
    -- CP-element group 232: 	230 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Sample/ack
      -- 
    ack_7650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3383_delayed_13_0_3474_inst_ack_0, ack => sendModule_CP_6819_elements(232)); -- 
    -- CP-element group 233:  transition  input  bypass  pipeline-parent 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	231 
    -- CP-element group 233: successors 
    -- CP-element group 233: 	358 
    -- CP-element group 233:  members (3) 
      -- CP-element group 233: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3476_Update/ack
      -- 
    ack_7655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3383_delayed_13_0_3474_inst_ack_1, ack => sendModule_CP_6819_elements(233)); -- 
    -- CP-element group 234:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	26 
    -- CP-element group 234: marked-predecessors 
    -- CP-element group 234: 	236 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (3) 
      -- CP-element group 234: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_sample_start_
      -- CP-element group 234: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Sample/$entry
      -- CP-element group 234: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Sample/rr
      -- 
    rr_7663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(234), ack => EQ_u3_u1_3486_inst_req_0); -- 
    sendModule_cp_element_group_234: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_234"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(236);
      gj_sendModule_cp_element_group_234 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(234), clk => clk, reset => reset); --
    end block;
    -- CP-element group 235:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: marked-predecessors 
    -- CP-element group 235: 	360 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	237 
    -- CP-element group 235:  members (3) 
      -- CP-element group 235: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_update_start_
      -- CP-element group 235: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Update/$entry
      -- CP-element group 235: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Update/cr
      -- 
    cr_7668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(235), ack => EQ_u3_u1_3486_inst_req_1); -- 
    sendModule_cp_element_group_235: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_235"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_235 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(235), clk => clk, reset => reset); --
    end block;
    -- CP-element group 236:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: successors 
    -- CP-element group 236: marked-successors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	22 
    -- CP-element group 236:  members (3) 
      -- CP-element group 236: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_sample_completed_
      -- CP-element group 236: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Sample/$exit
      -- CP-element group 236: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Sample/ra
      -- 
    ra_7664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 236_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3486_inst_ack_0, ack => sendModule_CP_6819_elements(236)); -- 
    -- CP-element group 237:  transition  input  bypass  pipeline-parent 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	235 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	358 
    -- CP-element group 237:  members (3) 
      -- CP-element group 237: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_update_completed_
      -- CP-element group 237: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Update/$exit
      -- CP-element group 237: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3486_Update/ca
      -- 
    ca_7669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3486_inst_ack_1, ack => sendModule_CP_6819_elements(237)); -- 
    -- CP-element group 238:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	157 
    -- CP-element group 238: marked-predecessors 
    -- CP-element group 238: 	240 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	240 
    -- CP-element group 238:  members (3) 
      -- CP-element group 238: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_sample_start_
      -- CP-element group 238: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Sample/$entry
      -- CP-element group 238: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Sample/req
      -- 
    req_7677_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7677_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(238), ack => W_output_data1_3391_delayed_13_0_3488_inst_req_0); -- 
    sendModule_cp_element_group_238: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_238"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(240);
      gj_sendModule_cp_element_group_238 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(238), clk => clk, reset => reset); --
    end block;
    -- CP-element group 239:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: marked-predecessors 
    -- CP-element group 239: 	360 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	241 
    -- CP-element group 239:  members (3) 
      -- CP-element group 239: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_update_start_
      -- CP-element group 239: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Update/$entry
      -- CP-element group 239: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Update/req
      -- 
    req_7682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(239), ack => W_output_data1_3391_delayed_13_0_3488_inst_req_1); -- 
    sendModule_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	238 
    -- CP-element group 240: successors 
    -- CP-element group 240: marked-successors 
    -- CP-element group 240: 	155 
    -- CP-element group 240: 	238 
    -- CP-element group 240:  members (3) 
      -- CP-element group 240: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_sample_completed_
      -- CP-element group 240: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Sample/$exit
      -- CP-element group 240: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Sample/ack
      -- 
    ack_7678_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 240_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3391_delayed_13_0_3488_inst_ack_0, ack => sendModule_CP_6819_elements(240)); -- 
    -- CP-element group 241:  transition  input  bypass  pipeline-parent 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	239 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	358 
    -- CP-element group 241:  members (3) 
      -- CP-element group 241: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_update_completed_
      -- CP-element group 241: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Update/$exit
      -- CP-element group 241: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3490_Update/ack
      -- 
    ack_7683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 241_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3391_delayed_13_0_3488_inst_ack_1, ack => sendModule_CP_6819_elements(241)); -- 
    -- CP-element group 242:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	26 
    -- CP-element group 242: marked-predecessors 
    -- CP-element group 242: 	244 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (3) 
      -- CP-element group 242: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_sample_start_
      -- CP-element group 242: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Sample/$entry
      -- CP-element group 242: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Sample/rr
      -- 
    rr_7691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(242), ack => EQ_u3_u1_3500_inst_req_0); -- 
    sendModule_cp_element_group_242: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_242"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(244);
      gj_sendModule_cp_element_group_242 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(242), clk => clk, reset => reset); --
    end block;
    -- CP-element group 243:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: marked-predecessors 
    -- CP-element group 243: 	360 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	245 
    -- CP-element group 243:  members (3) 
      -- CP-element group 243: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_update_start_
      -- CP-element group 243: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Update/$entry
      -- CP-element group 243: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Update/cr
      -- 
    cr_7696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(243), ack => EQ_u3_u1_3500_inst_req_1); -- 
    sendModule_cp_element_group_243: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_243"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_243 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(243), clk => clk, reset => reset); --
    end block;
    -- CP-element group 244:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: successors 
    -- CP-element group 244: marked-successors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	22 
    -- CP-element group 244:  members (3) 
      -- CP-element group 244: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_sample_completed_
      -- CP-element group 244: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Sample/$exit
      -- CP-element group 244: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Sample/ra
      -- 
    ra_7692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 244_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3500_inst_ack_0, ack => sendModule_CP_6819_elements(244)); -- 
    -- CP-element group 245:  transition  input  bypass  pipeline-parent 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	243 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	358 
    -- CP-element group 245:  members (3) 
      -- CP-element group 245: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_update_completed_
      -- CP-element group 245: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Update/$exit
      -- CP-element group 245: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3500_Update/ca
      -- 
    ca_7697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 245_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3500_inst_ack_1, ack => sendModule_CP_6819_elements(245)); -- 
    -- CP-element group 246:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	157 
    -- CP-element group 246: marked-predecessors 
    -- CP-element group 246: 	248 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (3) 
      -- CP-element group 246: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_sample_start_
      -- CP-element group 246: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Sample/$entry
      -- CP-element group 246: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Sample/req
      -- 
    req_7705_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7705_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(246), ack => W_output_data1_3399_delayed_13_0_3502_inst_req_0); -- 
    sendModule_cp_element_group_246: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_246"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(248);
      gj_sendModule_cp_element_group_246 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(246), clk => clk, reset => reset); --
    end block;
    -- CP-element group 247:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: marked-predecessors 
    -- CP-element group 247: 	360 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (3) 
      -- CP-element group 247: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_update_start_
      -- CP-element group 247: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Update/$entry
      -- CP-element group 247: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Update/req
      -- 
    req_7710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(247), ack => W_output_data1_3399_delayed_13_0_3502_inst_req_1); -- 
    sendModule_cp_element_group_247: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_247"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_247 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(247), clk => clk, reset => reset); --
    end block;
    -- CP-element group 248:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: marked-successors 
    -- CP-element group 248: 	155 
    -- CP-element group 248: 	246 
    -- CP-element group 248:  members (3) 
      -- CP-element group 248: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_sample_completed_
      -- CP-element group 248: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Sample/$exit
      -- CP-element group 248: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Sample/ack
      -- 
    ack_7706_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3399_delayed_13_0_3502_inst_ack_0, ack => sendModule_CP_6819_elements(248)); -- 
    -- CP-element group 249:  transition  input  bypass  pipeline-parent 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	358 
    -- CP-element group 249:  members (3) 
      -- CP-element group 249: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_update_completed_
      -- CP-element group 249: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Update/$exit
      -- CP-element group 249: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3504_Update/ack
      -- 
    ack_7711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 249_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3399_delayed_13_0_3502_inst_ack_1, ack => sendModule_CP_6819_elements(249)); -- 
    -- CP-element group 250:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	26 
    -- CP-element group 250: marked-predecessors 
    -- CP-element group 250: 	252 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (3) 
      -- CP-element group 250: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_sample_start_
      -- CP-element group 250: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Sample/$entry
      -- CP-element group 250: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Sample/rr
      -- 
    rr_7719_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7719_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(250), ack => EQ_u3_u1_3514_inst_req_0); -- 
    sendModule_cp_element_group_250: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_250"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(252);
      gj_sendModule_cp_element_group_250 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(250), clk => clk, reset => reset); --
    end block;
    -- CP-element group 251:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: marked-predecessors 
    -- CP-element group 251: 	360 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	253 
    -- CP-element group 251:  members (3) 
      -- CP-element group 251: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_update_start_
      -- CP-element group 251: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Update/$entry
      -- CP-element group 251: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Update/cr
      -- 
    cr_7724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(251), ack => EQ_u3_u1_3514_inst_req_1); -- 
    sendModule_cp_element_group_251: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_251"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_251 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(251), clk => clk, reset => reset); --
    end block;
    -- CP-element group 252:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: successors 
    -- CP-element group 252: marked-successors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	22 
    -- CP-element group 252:  members (3) 
      -- CP-element group 252: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_sample_completed_
      -- CP-element group 252: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Sample/$exit
      -- CP-element group 252: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Sample/ra
      -- 
    ra_7720_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 252_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3514_inst_ack_0, ack => sendModule_CP_6819_elements(252)); -- 
    -- CP-element group 253:  transition  input  bypass  pipeline-parent 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	251 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	358 
    -- CP-element group 253:  members (3) 
      -- CP-element group 253: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_update_completed_
      -- CP-element group 253: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Update/$exit
      -- CP-element group 253: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3514_Update/ca
      -- 
    ca_7725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3514_inst_ack_1, ack => sendModule_CP_6819_elements(253)); -- 
    -- CP-element group 254:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	157 
    -- CP-element group 254: marked-predecessors 
    -- CP-element group 254: 	256 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (3) 
      -- CP-element group 254: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_sample_start_
      -- CP-element group 254: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Sample/$entry
      -- CP-element group 254: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Sample/req
      -- 
    req_7733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(254), ack => W_output_data1_3407_delayed_13_0_3516_inst_req_0); -- 
    sendModule_cp_element_group_254: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_254"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(256);
      gj_sendModule_cp_element_group_254 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(254), clk => clk, reset => reset); --
    end block;
    -- CP-element group 255:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: marked-predecessors 
    -- CP-element group 255: 	360 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	257 
    -- CP-element group 255:  members (3) 
      -- CP-element group 255: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_update_start_
      -- CP-element group 255: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Update/$entry
      -- CP-element group 255: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Update/req
      -- 
    req_7738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(255), ack => W_output_data1_3407_delayed_13_0_3516_inst_req_1); -- 
    sendModule_cp_element_group_255: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_255"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_255 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(255), clk => clk, reset => reset); --
    end block;
    -- CP-element group 256:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: successors 
    -- CP-element group 256: marked-successors 
    -- CP-element group 256: 	155 
    -- CP-element group 256: 	254 
    -- CP-element group 256:  members (3) 
      -- CP-element group 256: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_sample_completed_
      -- CP-element group 256: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Sample/$exit
      -- CP-element group 256: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Sample/ack
      -- 
    ack_7734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 256_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3407_delayed_13_0_3516_inst_ack_0, ack => sendModule_CP_6819_elements(256)); -- 
    -- CP-element group 257:  transition  input  bypass  pipeline-parent 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	255 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	358 
    -- CP-element group 257:  members (3) 
      -- CP-element group 257: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_update_completed_
      -- CP-element group 257: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Update/$exit
      -- CP-element group 257: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3518_Update/ack
      -- 
    ack_7739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3407_delayed_13_0_3516_inst_ack_1, ack => sendModule_CP_6819_elements(257)); -- 
    -- CP-element group 258:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	26 
    -- CP-element group 258: marked-predecessors 
    -- CP-element group 258: 	260 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	260 
    -- CP-element group 258:  members (3) 
      -- CP-element group 258: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_sample_start_
      -- CP-element group 258: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Sample/$entry
      -- CP-element group 258: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Sample/rr
      -- 
    rr_7747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(258), ack => EQ_u3_u1_3528_inst_req_0); -- 
    sendModule_cp_element_group_258: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_258"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(260);
      gj_sendModule_cp_element_group_258 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(258), clk => clk, reset => reset); --
    end block;
    -- CP-element group 259:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: marked-predecessors 
    -- CP-element group 259: 	360 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	261 
    -- CP-element group 259:  members (3) 
      -- CP-element group 259: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_update_start_
      -- CP-element group 259: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Update/$entry
      -- CP-element group 259: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Update/cr
      -- 
    cr_7752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(259), ack => EQ_u3_u1_3528_inst_req_1); -- 
    sendModule_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: successors 
    -- CP-element group 260: marked-successors 
    -- CP-element group 260: 	258 
    -- CP-element group 260: 	22 
    -- CP-element group 260:  members (3) 
      -- CP-element group 260: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_sample_completed_
      -- CP-element group 260: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Sample/$exit
      -- CP-element group 260: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Sample/ra
      -- 
    ra_7748_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 260_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3528_inst_ack_0, ack => sendModule_CP_6819_elements(260)); -- 
    -- CP-element group 261:  transition  input  bypass  pipeline-parent 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	259 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	358 
    -- CP-element group 261:  members (3) 
      -- CP-element group 261: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_update_completed_
      -- CP-element group 261: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Update/$exit
      -- CP-element group 261: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3528_Update/ca
      -- 
    ca_7753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3528_inst_ack_1, ack => sendModule_CP_6819_elements(261)); -- 
    -- CP-element group 262:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	157 
    -- CP-element group 262: marked-predecessors 
    -- CP-element group 262: 	264 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (3) 
      -- CP-element group 262: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_sample_start_
      -- CP-element group 262: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Sample/$entry
      -- CP-element group 262: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Sample/req
      -- 
    req_7761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(262), ack => W_output_data1_3415_delayed_13_0_3530_inst_req_0); -- 
    sendModule_cp_element_group_262: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_262"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(264);
      gj_sendModule_cp_element_group_262 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(262), clk => clk, reset => reset); --
    end block;
    -- CP-element group 263:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: marked-predecessors 
    -- CP-element group 263: 	360 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	265 
    -- CP-element group 263:  members (3) 
      -- CP-element group 263: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_update_start_
      -- CP-element group 263: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Update/$entry
      -- CP-element group 263: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Update/req
      -- 
    req_7766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(263), ack => W_output_data1_3415_delayed_13_0_3530_inst_req_1); -- 
    sendModule_cp_element_group_263: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_263"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_263 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(263), clk => clk, reset => reset); --
    end block;
    -- CP-element group 264:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: successors 
    -- CP-element group 264: marked-successors 
    -- CP-element group 264: 	155 
    -- CP-element group 264: 	262 
    -- CP-element group 264:  members (3) 
      -- CP-element group 264: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_sample_completed_
      -- CP-element group 264: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Sample/$exit
      -- CP-element group 264: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Sample/ack
      -- 
    ack_7762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 264_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3415_delayed_13_0_3530_inst_ack_0, ack => sendModule_CP_6819_elements(264)); -- 
    -- CP-element group 265:  transition  input  bypass  pipeline-parent 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	263 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	358 
    -- CP-element group 265:  members (3) 
      -- CP-element group 265: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_update_completed_
      -- CP-element group 265: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Update/$exit
      -- CP-element group 265: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3532_Update/ack
      -- 
    ack_7767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 265_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3415_delayed_13_0_3530_inst_ack_1, ack => sendModule_CP_6819_elements(265)); -- 
    -- CP-element group 266:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	26 
    -- CP-element group 266: marked-predecessors 
    -- CP-element group 266: 	268 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	268 
    -- CP-element group 266:  members (3) 
      -- CP-element group 266: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_sample_start_
      -- CP-element group 266: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Sample/$entry
      -- CP-element group 266: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Sample/rr
      -- 
    rr_7775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(266), ack => EQ_u3_u1_3542_inst_req_0); -- 
    sendModule_cp_element_group_266: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_266"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(268);
      gj_sendModule_cp_element_group_266 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(266), clk => clk, reset => reset); --
    end block;
    -- CP-element group 267:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: marked-predecessors 
    -- CP-element group 267: 	360 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	269 
    -- CP-element group 267:  members (3) 
      -- CP-element group 267: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_update_start_
      -- CP-element group 267: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Update/cr
      -- 
    cr_7780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(267), ack => EQ_u3_u1_3542_inst_req_1); -- 
    sendModule_cp_element_group_267: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_267"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_267 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(267), clk => clk, reset => reset); --
    end block;
    -- CP-element group 268:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: successors 
    -- CP-element group 268: marked-successors 
    -- CP-element group 268: 	266 
    -- CP-element group 268: 	22 
    -- CP-element group 268:  members (3) 
      -- CP-element group 268: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_sample_completed_
      -- CP-element group 268: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Sample/$exit
      -- CP-element group 268: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Sample/ra
      -- 
    ra_7776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 268_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3542_inst_ack_0, ack => sendModule_CP_6819_elements(268)); -- 
    -- CP-element group 269:  transition  input  bypass  pipeline-parent 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	267 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	358 
    -- CP-element group 269:  members (3) 
      -- CP-element group 269: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_update_completed_
      -- CP-element group 269: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Update/$exit
      -- CP-element group 269: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3542_Update/ca
      -- 
    ca_7781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 269_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3542_inst_ack_1, ack => sendModule_CP_6819_elements(269)); -- 
    -- CP-element group 270:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	157 
    -- CP-element group 270: marked-predecessors 
    -- CP-element group 270: 	272 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (3) 
      -- CP-element group 270: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_sample_start_
      -- CP-element group 270: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Sample/$entry
      -- CP-element group 270: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Sample/req
      -- 
    req_7789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(270), ack => W_output_data1_3423_delayed_13_0_3544_inst_req_0); -- 
    sendModule_cp_element_group_270: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_270"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(272);
      gj_sendModule_cp_element_group_270 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(270), clk => clk, reset => reset); --
    end block;
    -- CP-element group 271:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: marked-predecessors 
    -- CP-element group 271: 	360 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	273 
    -- CP-element group 271:  members (3) 
      -- CP-element group 271: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_update_start_
      -- CP-element group 271: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Update/$entry
      -- CP-element group 271: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Update/req
      -- 
    req_7794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(271), ack => W_output_data1_3423_delayed_13_0_3544_inst_req_1); -- 
    sendModule_cp_element_group_271: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_271"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_271 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(271), clk => clk, reset => reset); --
    end block;
    -- CP-element group 272:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: successors 
    -- CP-element group 272: marked-successors 
    -- CP-element group 272: 	155 
    -- CP-element group 272: 	270 
    -- CP-element group 272:  members (3) 
      -- CP-element group 272: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_sample_completed_
      -- CP-element group 272: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Sample/$exit
      -- CP-element group 272: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Sample/ack
      -- 
    ack_7790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 272_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3423_delayed_13_0_3544_inst_ack_0, ack => sendModule_CP_6819_elements(272)); -- 
    -- CP-element group 273:  transition  input  bypass  pipeline-parent 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	271 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	358 
    -- CP-element group 273:  members (3) 
      -- CP-element group 273: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_update_completed_
      -- CP-element group 273: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Update/$exit
      -- CP-element group 273: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3546_Update/ack
      -- 
    ack_7795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 273_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3423_delayed_13_0_3544_inst_ack_1, ack => sendModule_CP_6819_elements(273)); -- 
    -- CP-element group 274:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	26 
    -- CP-element group 274: marked-predecessors 
    -- CP-element group 274: 	276 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (3) 
      -- CP-element group 274: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Sample/rr
      -- CP-element group 274: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Sample/$entry
      -- CP-element group 274: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_sample_start_
      -- 
    rr_7803_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7803_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(274), ack => EQ_u3_u1_3556_inst_req_0); -- 
    sendModule_cp_element_group_274: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_274"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(276);
      gj_sendModule_cp_element_group_274 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(274), clk => clk, reset => reset); --
    end block;
    -- CP-element group 275:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: marked-predecessors 
    -- CP-element group 275: 	360 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	277 
    -- CP-element group 275:  members (3) 
      -- CP-element group 275: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Update/cr
      -- CP-element group 275: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Update/$entry
      -- CP-element group 275: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_update_start_
      -- 
    cr_7808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(275), ack => EQ_u3_u1_3556_inst_req_1); -- 
    sendModule_cp_element_group_275: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_275"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_275 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(275), clk => clk, reset => reset); --
    end block;
    -- CP-element group 276:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: successors 
    -- CP-element group 276: marked-successors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	22 
    -- CP-element group 276:  members (3) 
      -- CP-element group 276: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Sample/ra
      -- CP-element group 276: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Sample/$exit
      -- CP-element group 276: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_sample_completed_
      -- 
    ra_7804_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 276_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3556_inst_ack_0, ack => sendModule_CP_6819_elements(276)); -- 
    -- CP-element group 277:  transition  input  bypass  pipeline-parent 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	275 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	358 
    -- CP-element group 277:  members (3) 
      -- CP-element group 277: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Update/ca
      -- CP-element group 277: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_Update/$exit
      -- CP-element group 277: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3556_update_completed_
      -- 
    ca_7809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3556_inst_ack_1, ack => sendModule_CP_6819_elements(277)); -- 
    -- CP-element group 278:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	157 
    -- CP-element group 278: marked-predecessors 
    -- CP-element group 278: 	280 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	280 
    -- CP-element group 278:  members (3) 
      -- CP-element group 278: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Sample/req
      -- CP-element group 278: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Sample/$entry
      -- CP-element group 278: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_sample_start_
      -- 
    req_7817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(278), ack => W_output_data1_3431_delayed_13_0_3558_inst_req_0); -- 
    sendModule_cp_element_group_278: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_278"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(280);
      gj_sendModule_cp_element_group_278 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(278), clk => clk, reset => reset); --
    end block;
    -- CP-element group 279:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: marked-predecessors 
    -- CP-element group 279: 	360 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	281 
    -- CP-element group 279:  members (3) 
      -- CP-element group 279: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Update/$entry
      -- CP-element group 279: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_update_start_
      -- CP-element group 279: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Update/req
      -- 
    req_7822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(279), ack => W_output_data1_3431_delayed_13_0_3558_inst_req_1); -- 
    sendModule_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	278 
    -- CP-element group 280: successors 
    -- CP-element group 280: marked-successors 
    -- CP-element group 280: 	155 
    -- CP-element group 280: 	278 
    -- CP-element group 280:  members (3) 
      -- CP-element group 280: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Sample/ack
      -- CP-element group 280: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Sample/$exit
      -- CP-element group 280: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_sample_completed_
      -- 
    ack_7818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 280_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3431_delayed_13_0_3558_inst_ack_0, ack => sendModule_CP_6819_elements(280)); -- 
    -- CP-element group 281:  transition  input  bypass  pipeline-parent 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	279 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	358 
    -- CP-element group 281:  members (3) 
      -- CP-element group 281: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Update/$exit
      -- CP-element group 281: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_Update/ack
      -- CP-element group 281: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3560_update_completed_
      -- 
    ack_7823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 281_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3431_delayed_13_0_3558_inst_ack_1, ack => sendModule_CP_6819_elements(281)); -- 
    -- CP-element group 282:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	26 
    -- CP-element group 282: marked-predecessors 
    -- CP-element group 282: 	284 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (3) 
      -- CP-element group 282: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Sample/rr
      -- CP-element group 282: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Sample/$entry
      -- CP-element group 282: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_sample_start_
      -- 
    rr_7831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(282), ack => EQ_u3_u1_3570_inst_req_0); -- 
    sendModule_cp_element_group_282: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_282"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(26) & sendModule_CP_6819_elements(284);
      gj_sendModule_cp_element_group_282 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(282), clk => clk, reset => reset); --
    end block;
    -- CP-element group 283:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: marked-predecessors 
    -- CP-element group 283: 	360 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	285 
    -- CP-element group 283:  members (3) 
      -- CP-element group 283: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Update/$entry
      -- CP-element group 283: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_update_start_
      -- CP-element group 283: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Update/cr
      -- 
    cr_7836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(283), ack => EQ_u3_u1_3570_inst_req_1); -- 
    sendModule_cp_element_group_283: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_283"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_283 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(283), clk => clk, reset => reset); --
    end block;
    -- CP-element group 284:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: successors 
    -- CP-element group 284: marked-successors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	22 
    -- CP-element group 284:  members (3) 
      -- CP-element group 284: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Sample/ra
      -- CP-element group 284: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Sample/$exit
      -- CP-element group 284: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_sample_completed_
      -- 
    ra_7832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 284_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3570_inst_ack_0, ack => sendModule_CP_6819_elements(284)); -- 
    -- CP-element group 285:  transition  input  bypass  pipeline-parent 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	283 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	358 
    -- CP-element group 285:  members (3) 
      -- CP-element group 285: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Update/$exit
      -- CP-element group 285: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_update_completed_
      -- CP-element group 285: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3570_Update/ca
      -- 
    ca_7837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3570_inst_ack_1, ack => sendModule_CP_6819_elements(285)); -- 
    -- CP-element group 286:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	157 
    -- CP-element group 286: marked-predecessors 
    -- CP-element group 286: 	288 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	288 
    -- CP-element group 286:  members (3) 
      -- CP-element group 286: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Sample/req
      -- CP-element group 286: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Sample/$entry
      -- CP-element group 286: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_sample_start_
      -- 
    req_7845_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7845_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(286), ack => W_output_data1_3439_delayed_13_0_3572_inst_req_0); -- 
    sendModule_cp_element_group_286: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_286"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(157) & sendModule_CP_6819_elements(288);
      gj_sendModule_cp_element_group_286 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(286), clk => clk, reset => reset); --
    end block;
    -- CP-element group 287:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: marked-predecessors 
    -- CP-element group 287: 	360 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	289 
    -- CP-element group 287:  members (3) 
      -- CP-element group 287: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Update/req
      -- CP-element group 287: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Update/$entry
      -- CP-element group 287: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_update_start_
      -- 
    req_7850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(287), ack => W_output_data1_3439_delayed_13_0_3572_inst_req_1); -- 
    sendModule_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	286 
    -- CP-element group 288: successors 
    -- CP-element group 288: marked-successors 
    -- CP-element group 288: 	155 
    -- CP-element group 288: 	286 
    -- CP-element group 288:  members (3) 
      -- CP-element group 288: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Sample/ack
      -- CP-element group 288: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Sample/$exit
      -- CP-element group 288: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_sample_completed_
      -- 
    ack_7846_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3439_delayed_13_0_3572_inst_ack_0, ack => sendModule_CP_6819_elements(288)); -- 
    -- CP-element group 289:  transition  input  bypass  pipeline-parent 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	287 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	358 
    -- CP-element group 289:  members (3) 
      -- CP-element group 289: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Update/ack
      -- CP-element group 289: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_Update/$exit
      -- CP-element group 289: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3574_update_completed_
      -- 
    ack_7851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 289_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data1_3439_delayed_13_0_3572_inst_ack_1, ack => sendModule_CP_6819_elements(289)); -- 
    -- CP-element group 290:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	43 
    -- CP-element group 290: marked-predecessors 
    -- CP-element group 290: 	292 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	292 
    -- CP-element group 290:  members (3) 
      -- CP-element group 290: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Sample/$entry
      -- CP-element group 290: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Sample/rr
      -- CP-element group 290: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_sample_start_
      -- 
    rr_7859_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7859_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(290), ack => EQ_u3_u1_3584_inst_req_0); -- 
    sendModule_cp_element_group_290: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_290"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(292);
      gj_sendModule_cp_element_group_290 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(290), clk => clk, reset => reset); --
    end block;
    -- CP-element group 291:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: marked-predecessors 
    -- CP-element group 291: 	372 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (3) 
      -- CP-element group 291: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Update/$entry
      -- CP-element group 291: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_update_start_
      -- CP-element group 291: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Update/cr
      -- 
    cr_7864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(291), ack => EQ_u3_u1_3584_inst_req_1); -- 
    sendModule_cp_element_group_291: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_291"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_291 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(291), clk => clk, reset => reset); --
    end block;
    -- CP-element group 292:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: successors 
    -- CP-element group 292: marked-successors 
    -- CP-element group 292: 	290 
    -- CP-element group 292: 	41 
    -- CP-element group 292:  members (3) 
      -- CP-element group 292: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Sample/$exit
      -- CP-element group 292: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Sample/ra
      -- CP-element group 292: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_sample_completed_
      -- 
    ra_7860_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3584_inst_ack_0, ack => sendModule_CP_6819_elements(292)); -- 
    -- CP-element group 293:  transition  input  bypass  pipeline-parent 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	370 
    -- CP-element group 293:  members (3) 
      -- CP-element group 293: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Update/$exit
      -- CP-element group 293: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_update_completed_
      -- CP-element group 293: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3584_Update/ca
      -- 
    ca_7865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 293_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3584_inst_ack_1, ack => sendModule_CP_6819_elements(293)); -- 
    -- CP-element group 294:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	161 
    -- CP-element group 294: marked-predecessors 
    -- CP-element group 294: 	296 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	296 
    -- CP-element group 294:  members (3) 
      -- CP-element group 294: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Sample/req
      -- CP-element group 294: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Sample/$entry
      -- CP-element group 294: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_sample_start_
      -- 
    req_7873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(294), ack => W_output_data2_3447_delayed_13_0_3586_inst_req_0); -- 
    sendModule_cp_element_group_294: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_294"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(296);
      gj_sendModule_cp_element_group_294 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(294), clk => clk, reset => reset); --
    end block;
    -- CP-element group 295:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: marked-predecessors 
    -- CP-element group 295: 	372 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	297 
    -- CP-element group 295:  members (3) 
      -- CP-element group 295: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Update/req
      -- CP-element group 295: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_update_start_
      -- 
    req_7878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(295), ack => W_output_data2_3447_delayed_13_0_3586_inst_req_1); -- 
    sendModule_cp_element_group_295: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_295"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_295 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(295), clk => clk, reset => reset); --
    end block;
    -- CP-element group 296:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	294 
    -- CP-element group 296: successors 
    -- CP-element group 296: marked-successors 
    -- CP-element group 296: 	159 
    -- CP-element group 296: 	294 
    -- CP-element group 296:  members (3) 
      -- CP-element group 296: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Sample/ack
      -- CP-element group 296: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Sample/$exit
      -- CP-element group 296: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_sample_completed_
      -- 
    ack_7874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 296_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3447_delayed_13_0_3586_inst_ack_0, ack => sendModule_CP_6819_elements(296)); -- 
    -- CP-element group 297:  transition  input  bypass  pipeline-parent 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	295 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	370 
    -- CP-element group 297:  members (3) 
      -- CP-element group 297: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Update/ack
      -- CP-element group 297: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_Update/$exit
      -- CP-element group 297: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3588_update_completed_
      -- 
    ack_7879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3447_delayed_13_0_3586_inst_ack_1, ack => sendModule_CP_6819_elements(297)); -- 
    -- CP-element group 298:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	43 
    -- CP-element group 298: marked-predecessors 
    -- CP-element group 298: 	300 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	300 
    -- CP-element group 298:  members (3) 
      -- CP-element group 298: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Sample/rr
      -- CP-element group 298: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Sample/$entry
      -- CP-element group 298: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_sample_start_
      -- 
    rr_7887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(298), ack => EQ_u3_u1_3598_inst_req_0); -- 
    sendModule_cp_element_group_298: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_298"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(300);
      gj_sendModule_cp_element_group_298 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(298), clk => clk, reset => reset); --
    end block;
    -- CP-element group 299:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: marked-predecessors 
    -- CP-element group 299: 	372 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	301 
    -- CP-element group 299:  members (3) 
      -- CP-element group 299: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Update/cr
      -- CP-element group 299: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Update/$entry
      -- CP-element group 299: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_update_start_
      -- 
    cr_7892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(299), ack => EQ_u3_u1_3598_inst_req_1); -- 
    sendModule_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: successors 
    -- CP-element group 300: marked-successors 
    -- CP-element group 300: 	298 
    -- CP-element group 300: 	41 
    -- CP-element group 300:  members (3) 
      -- CP-element group 300: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Sample/ra
      -- CP-element group 300: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Sample/$exit
      -- CP-element group 300: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_sample_completed_
      -- 
    ra_7888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 300_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3598_inst_ack_0, ack => sendModule_CP_6819_elements(300)); -- 
    -- CP-element group 301:  transition  input  bypass  pipeline-parent 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	299 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	370 
    -- CP-element group 301:  members (3) 
      -- CP-element group 301: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Update/ca
      -- CP-element group 301: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_Update/$exit
      -- CP-element group 301: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3598_update_completed_
      -- 
    ca_7893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3598_inst_ack_1, ack => sendModule_CP_6819_elements(301)); -- 
    -- CP-element group 302:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	161 
    -- CP-element group 302: marked-predecessors 
    -- CP-element group 302: 	304 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	304 
    -- CP-element group 302:  members (3) 
      -- CP-element group 302: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Sample/$entry
      -- CP-element group 302: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Sample/req
      -- CP-element group 302: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_sample_start_
      -- 
    req_7901_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7901_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(302), ack => W_output_data2_3455_delayed_13_0_3600_inst_req_0); -- 
    sendModule_cp_element_group_302: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_302"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(304);
      gj_sendModule_cp_element_group_302 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(302), clk => clk, reset => reset); --
    end block;
    -- CP-element group 303:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: marked-predecessors 
    -- CP-element group 303: 	372 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	305 
    -- CP-element group 303:  members (3) 
      -- CP-element group 303: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Update/req
      -- CP-element group 303: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_update_start_
      -- 
    req_7906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(303), ack => W_output_data2_3455_delayed_13_0_3600_inst_req_1); -- 
    sendModule_cp_element_group_303: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_303"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_303 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(303), clk => clk, reset => reset); --
    end block;
    -- CP-element group 304:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	302 
    -- CP-element group 304: successors 
    -- CP-element group 304: marked-successors 
    -- CP-element group 304: 	159 
    -- CP-element group 304: 	302 
    -- CP-element group 304:  members (3) 
      -- CP-element group 304: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Sample/ack
      -- CP-element group 304: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Sample/$exit
      -- CP-element group 304: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_sample_completed_
      -- 
    ack_7902_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 304_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3455_delayed_13_0_3600_inst_ack_0, ack => sendModule_CP_6819_elements(304)); -- 
    -- CP-element group 305:  transition  input  bypass  pipeline-parent 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	303 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	370 
    -- CP-element group 305:  members (3) 
      -- CP-element group 305: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Update/$exit
      -- CP-element group 305: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_Update/ack
      -- CP-element group 305: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3602_update_completed_
      -- 
    ack_7907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3455_delayed_13_0_3600_inst_ack_1, ack => sendModule_CP_6819_elements(305)); -- 
    -- CP-element group 306:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	43 
    -- CP-element group 306: marked-predecessors 
    -- CP-element group 306: 	308 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	308 
    -- CP-element group 306:  members (3) 
      -- CP-element group 306: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_sample_start_
      -- CP-element group 306: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Sample/$entry
      -- CP-element group 306: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Sample/rr
      -- 
    rr_7915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(306), ack => EQ_u3_u1_3612_inst_req_0); -- 
    sendModule_cp_element_group_306: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_306"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(308);
      gj_sendModule_cp_element_group_306 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(306), clk => clk, reset => reset); --
    end block;
    -- CP-element group 307:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: marked-predecessors 
    -- CP-element group 307: 	372 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	309 
    -- CP-element group 307:  members (3) 
      -- CP-element group 307: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_update_start_
      -- CP-element group 307: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Update/cr
      -- CP-element group 307: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Update/$entry
      -- 
    cr_7920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(307), ack => EQ_u3_u1_3612_inst_req_1); -- 
    sendModule_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: successors 
    -- CP-element group 308: marked-successors 
    -- CP-element group 308: 	306 
    -- CP-element group 308: 	41 
    -- CP-element group 308:  members (3) 
      -- CP-element group 308: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_sample_completed_
      -- CP-element group 308: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Sample/ra
      -- CP-element group 308: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Sample/$exit
      -- 
    ra_7916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 308_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3612_inst_ack_0, ack => sendModule_CP_6819_elements(308)); -- 
    -- CP-element group 309:  transition  input  bypass  pipeline-parent 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	307 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	370 
    -- CP-element group 309:  members (3) 
      -- CP-element group 309: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_update_completed_
      -- CP-element group 309: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Update/ca
      -- CP-element group 309: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3612_Update/$exit
      -- 
    ca_7921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3612_inst_ack_1, ack => sendModule_CP_6819_elements(309)); -- 
    -- CP-element group 310:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	161 
    -- CP-element group 310: marked-predecessors 
    -- CP-element group 310: 	312 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	312 
    -- CP-element group 310:  members (3) 
      -- CP-element group 310: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Sample/req
      -- CP-element group 310: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_sample_start_
      -- 
    req_7929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(310), ack => W_output_data2_3463_delayed_13_0_3614_inst_req_0); -- 
    sendModule_cp_element_group_310: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_310"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(312);
      gj_sendModule_cp_element_group_310 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(310), clk => clk, reset => reset); --
    end block;
    -- CP-element group 311:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 311: predecessors 
    -- CP-element group 311: marked-predecessors 
    -- CP-element group 311: 	372 
    -- CP-element group 311: successors 
    -- CP-element group 311: 	313 
    -- CP-element group 311:  members (3) 
      -- CP-element group 311: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Update/req
      -- CP-element group 311: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Update/$entry
      -- CP-element group 311: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_update_start_
      -- 
    req_7934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(311), ack => W_output_data2_3463_delayed_13_0_3614_inst_req_1); -- 
    sendModule_cp_element_group_311: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_311"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_311 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(311), clk => clk, reset => reset); --
    end block;
    -- CP-element group 312:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 312: predecessors 
    -- CP-element group 312: 	310 
    -- CP-element group 312: successors 
    -- CP-element group 312: marked-successors 
    -- CP-element group 312: 	159 
    -- CP-element group 312: 	310 
    -- CP-element group 312:  members (3) 
      -- CP-element group 312: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Sample/ack
      -- CP-element group 312: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Sample/$exit
      -- CP-element group 312: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_sample_completed_
      -- 
    ack_7930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 312_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3463_delayed_13_0_3614_inst_ack_0, ack => sendModule_CP_6819_elements(312)); -- 
    -- CP-element group 313:  transition  input  bypass  pipeline-parent 
    -- CP-element group 313: predecessors 
    -- CP-element group 313: 	311 
    -- CP-element group 313: successors 
    -- CP-element group 313: 	370 
    -- CP-element group 313:  members (3) 
      -- CP-element group 313: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Update/ack
      -- CP-element group 313: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_Update/$exit
      -- CP-element group 313: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3616_update_completed_
      -- 
    ack_7935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 313_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3463_delayed_13_0_3614_inst_ack_1, ack => sendModule_CP_6819_elements(313)); -- 
    -- CP-element group 314:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 314: predecessors 
    -- CP-element group 314: 	43 
    -- CP-element group 314: marked-predecessors 
    -- CP-element group 314: 	316 
    -- CP-element group 314: successors 
    -- CP-element group 314: 	316 
    -- CP-element group 314:  members (3) 
      -- CP-element group 314: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Sample/rr
      -- CP-element group 314: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Sample/$entry
      -- CP-element group 314: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_sample_start_
      -- 
    rr_7943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(314), ack => EQ_u3_u1_3626_inst_req_0); -- 
    sendModule_cp_element_group_314: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_314"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(316);
      gj_sendModule_cp_element_group_314 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(314), clk => clk, reset => reset); --
    end block;
    -- CP-element group 315:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 315: predecessors 
    -- CP-element group 315: marked-predecessors 
    -- CP-element group 315: 	372 
    -- CP-element group 315: successors 
    -- CP-element group 315: 	317 
    -- CP-element group 315:  members (3) 
      -- CP-element group 315: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Update/cr
      -- CP-element group 315: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Update/$entry
      -- CP-element group 315: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_update_start_
      -- 
    cr_7948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(315), ack => EQ_u3_u1_3626_inst_req_1); -- 
    sendModule_cp_element_group_315: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_315"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_315 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(315), clk => clk, reset => reset); --
    end block;
    -- CP-element group 316:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 316: predecessors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: successors 
    -- CP-element group 316: marked-successors 
    -- CP-element group 316: 	314 
    -- CP-element group 316: 	41 
    -- CP-element group 316:  members (3) 
      -- CP-element group 316: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Sample/ra
      -- CP-element group 316: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Sample/$exit
      -- CP-element group 316: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_sample_completed_
      -- 
    ra_7944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 316_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3626_inst_ack_0, ack => sendModule_CP_6819_elements(316)); -- 
    -- CP-element group 317:  transition  input  bypass  pipeline-parent 
    -- CP-element group 317: predecessors 
    -- CP-element group 317: 	315 
    -- CP-element group 317: successors 
    -- CP-element group 317: 	370 
    -- CP-element group 317:  members (3) 
      -- CP-element group 317: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Update/ca
      -- CP-element group 317: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_Update/$exit
      -- CP-element group 317: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3626_update_completed_
      -- 
    ca_7949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 317_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3626_inst_ack_1, ack => sendModule_CP_6819_elements(317)); -- 
    -- CP-element group 318:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 318: predecessors 
    -- CP-element group 318: 	161 
    -- CP-element group 318: marked-predecessors 
    -- CP-element group 318: 	320 
    -- CP-element group 318: successors 
    -- CP-element group 318: 	320 
    -- CP-element group 318:  members (3) 
      -- CP-element group 318: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Sample/$entry
      -- CP-element group 318: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_sample_start_
      -- CP-element group 318: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Sample/req
      -- 
    req_7957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(318), ack => W_output_data2_3471_delayed_13_0_3628_inst_req_0); -- 
    sendModule_cp_element_group_318: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_318"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(320);
      gj_sendModule_cp_element_group_318 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(318), clk => clk, reset => reset); --
    end block;
    -- CP-element group 319:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 319: predecessors 
    -- CP-element group 319: marked-predecessors 
    -- CP-element group 319: 	372 
    -- CP-element group 319: successors 
    -- CP-element group 319: 	321 
    -- CP-element group 319:  members (3) 
      -- CP-element group 319: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_update_start_
      -- CP-element group 319: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Update/req
      -- CP-element group 319: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Update/$entry
      -- 
    req_7962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(319), ack => W_output_data2_3471_delayed_13_0_3628_inst_req_1); -- 
    sendModule_cp_element_group_319: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_319"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_319 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(319), clk => clk, reset => reset); --
    end block;
    -- CP-element group 320:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 320: predecessors 
    -- CP-element group 320: 	318 
    -- CP-element group 320: successors 
    -- CP-element group 320: marked-successors 
    -- CP-element group 320: 	159 
    -- CP-element group 320: 	318 
    -- CP-element group 320:  members (3) 
      -- CP-element group 320: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Sample/$exit
      -- CP-element group 320: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_sample_completed_
      -- CP-element group 320: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Sample/ack
      -- 
    ack_7958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 320_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3471_delayed_13_0_3628_inst_ack_0, ack => sendModule_CP_6819_elements(320)); -- 
    -- CP-element group 321:  transition  input  bypass  pipeline-parent 
    -- CP-element group 321: predecessors 
    -- CP-element group 321: 	319 
    -- CP-element group 321: successors 
    -- CP-element group 321: 	370 
    -- CP-element group 321:  members (3) 
      -- CP-element group 321: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_update_completed_
      -- CP-element group 321: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Update/ack
      -- CP-element group 321: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3630_Update/$exit
      -- 
    ack_7963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 321_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3471_delayed_13_0_3628_inst_ack_1, ack => sendModule_CP_6819_elements(321)); -- 
    -- CP-element group 322:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 322: predecessors 
    -- CP-element group 322: 	43 
    -- CP-element group 322: marked-predecessors 
    -- CP-element group 322: 	324 
    -- CP-element group 322: successors 
    -- CP-element group 322: 	324 
    -- CP-element group 322:  members (3) 
      -- CP-element group 322: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Sample/rr
      -- CP-element group 322: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Sample/$entry
      -- CP-element group 322: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_sample_start_
      -- 
    rr_7971_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7971_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(322), ack => EQ_u3_u1_3640_inst_req_0); -- 
    sendModule_cp_element_group_322: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_322"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(324);
      gj_sendModule_cp_element_group_322 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(322), clk => clk, reset => reset); --
    end block;
    -- CP-element group 323:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 323: predecessors 
    -- CP-element group 323: marked-predecessors 
    -- CP-element group 323: 	372 
    -- CP-element group 323: successors 
    -- CP-element group 323: 	325 
    -- CP-element group 323:  members (3) 
      -- CP-element group 323: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Update/cr
      -- CP-element group 323: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Update/$entry
      -- CP-element group 323: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_update_start_
      -- 
    cr_7976_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7976_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(323), ack => EQ_u3_u1_3640_inst_req_1); -- 
    sendModule_cp_element_group_323: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_323"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_323 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(323), clk => clk, reset => reset); --
    end block;
    -- CP-element group 324:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 324: predecessors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: successors 
    -- CP-element group 324: marked-successors 
    -- CP-element group 324: 	322 
    -- CP-element group 324: 	41 
    -- CP-element group 324:  members (3) 
      -- CP-element group 324: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Sample/ra
      -- CP-element group 324: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Sample/$exit
      -- CP-element group 324: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_sample_completed_
      -- 
    ra_7972_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 324_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3640_inst_ack_0, ack => sendModule_CP_6819_elements(324)); -- 
    -- CP-element group 325:  transition  input  bypass  pipeline-parent 
    -- CP-element group 325: predecessors 
    -- CP-element group 325: 	323 
    -- CP-element group 325: successors 
    -- CP-element group 325: 	370 
    -- CP-element group 325:  members (3) 
      -- CP-element group 325: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Update/ca
      -- CP-element group 325: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_Update/$exit
      -- CP-element group 325: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3640_update_completed_
      -- 
    ca_7977_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 325_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3640_inst_ack_1, ack => sendModule_CP_6819_elements(325)); -- 
    -- CP-element group 326:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 326: predecessors 
    -- CP-element group 326: 	161 
    -- CP-element group 326: marked-predecessors 
    -- CP-element group 326: 	328 
    -- CP-element group 326: successors 
    -- CP-element group 326: 	328 
    -- CP-element group 326:  members (3) 
      -- CP-element group 326: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Sample/$entry
      -- CP-element group 326: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Sample/req
      -- CP-element group 326: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_sample_start_
      -- 
    req_7985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(326), ack => W_output_data2_3479_delayed_13_0_3642_inst_req_0); -- 
    sendModule_cp_element_group_326: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_326"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(328);
      gj_sendModule_cp_element_group_326 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(326), clk => clk, reset => reset); --
    end block;
    -- CP-element group 327:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 327: predecessors 
    -- CP-element group 327: marked-predecessors 
    -- CP-element group 327: 	372 
    -- CP-element group 327: successors 
    -- CP-element group 327: 	329 
    -- CP-element group 327:  members (3) 
      -- CP-element group 327: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Update/$entry
      -- CP-element group 327: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Update/req
      -- CP-element group 327: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_update_start_
      -- 
    req_7990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(327), ack => W_output_data2_3479_delayed_13_0_3642_inst_req_1); -- 
    sendModule_cp_element_group_327: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_327"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_327 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(327), clk => clk, reset => reset); --
    end block;
    -- CP-element group 328:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 328: predecessors 
    -- CP-element group 328: 	326 
    -- CP-element group 328: successors 
    -- CP-element group 328: marked-successors 
    -- CP-element group 328: 	159 
    -- CP-element group 328: 	326 
    -- CP-element group 328:  members (3) 
      -- CP-element group 328: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Sample/$exit
      -- CP-element group 328: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Sample/ack
      -- CP-element group 328: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_sample_completed_
      -- 
    ack_7986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 328_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3479_delayed_13_0_3642_inst_ack_0, ack => sendModule_CP_6819_elements(328)); -- 
    -- CP-element group 329:  transition  input  bypass  pipeline-parent 
    -- CP-element group 329: predecessors 
    -- CP-element group 329: 	327 
    -- CP-element group 329: successors 
    -- CP-element group 329: 	370 
    -- CP-element group 329:  members (3) 
      -- CP-element group 329: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Update/$exit
      -- CP-element group 329: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_Update/ack
      -- CP-element group 329: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3644_update_completed_
      -- 
    ack_7991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 329_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3479_delayed_13_0_3642_inst_ack_1, ack => sendModule_CP_6819_elements(329)); -- 
    -- CP-element group 330:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 330: predecessors 
    -- CP-element group 330: 	43 
    -- CP-element group 330: marked-predecessors 
    -- CP-element group 330: 	332 
    -- CP-element group 330: successors 
    -- CP-element group 330: 	332 
    -- CP-element group 330:  members (3) 
      -- CP-element group 330: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_sample_start_
      -- CP-element group 330: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Sample/rr
      -- CP-element group 330: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Sample/$entry
      -- 
    rr_7999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(330), ack => EQ_u3_u1_3654_inst_req_0); -- 
    sendModule_cp_element_group_330: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_330"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(332);
      gj_sendModule_cp_element_group_330 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(330), clk => clk, reset => reset); --
    end block;
    -- CP-element group 331:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 331: predecessors 
    -- CP-element group 331: marked-predecessors 
    -- CP-element group 331: 	372 
    -- CP-element group 331: successors 
    -- CP-element group 331: 	333 
    -- CP-element group 331:  members (3) 
      -- CP-element group 331: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Update/cr
      -- CP-element group 331: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Update/$entry
      -- CP-element group 331: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_update_start_
      -- 
    cr_8004_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8004_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(331), ack => EQ_u3_u1_3654_inst_req_1); -- 
    sendModule_cp_element_group_331: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_331"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_331 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(331), clk => clk, reset => reset); --
    end block;
    -- CP-element group 332:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 332: predecessors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: successors 
    -- CP-element group 332: marked-successors 
    -- CP-element group 332: 	330 
    -- CP-element group 332: 	41 
    -- CP-element group 332:  members (3) 
      -- CP-element group 332: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Sample/ra
      -- CP-element group 332: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Sample/$exit
      -- CP-element group 332: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_sample_completed_
      -- 
    ra_8000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 332_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3654_inst_ack_0, ack => sendModule_CP_6819_elements(332)); -- 
    -- CP-element group 333:  transition  input  bypass  pipeline-parent 
    -- CP-element group 333: predecessors 
    -- CP-element group 333: 	331 
    -- CP-element group 333: successors 
    -- CP-element group 333: 	370 
    -- CP-element group 333:  members (3) 
      -- CP-element group 333: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Update/ca
      -- CP-element group 333: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_Update/$exit
      -- CP-element group 333: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3654_update_completed_
      -- 
    ca_8005_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 333_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3654_inst_ack_1, ack => sendModule_CP_6819_elements(333)); -- 
    -- CP-element group 334:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 334: predecessors 
    -- CP-element group 334: 	161 
    -- CP-element group 334: marked-predecessors 
    -- CP-element group 334: 	336 
    -- CP-element group 334: successors 
    -- CP-element group 334: 	336 
    -- CP-element group 334:  members (3) 
      -- CP-element group 334: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_sample_start_
      -- CP-element group 334: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Sample/req
      -- CP-element group 334: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Sample/$entry
      -- 
    req_8013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(334), ack => W_output_data2_3487_delayed_13_0_3656_inst_req_0); -- 
    sendModule_cp_element_group_334: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_334"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(336);
      gj_sendModule_cp_element_group_334 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(334), clk => clk, reset => reset); --
    end block;
    -- CP-element group 335:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 335: predecessors 
    -- CP-element group 335: marked-predecessors 
    -- CP-element group 335: 	372 
    -- CP-element group 335: successors 
    -- CP-element group 335: 	337 
    -- CP-element group 335:  members (3) 
      -- CP-element group 335: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_update_start_
      -- CP-element group 335: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Update/req
      -- CP-element group 335: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Update/$entry
      -- 
    req_8018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(335), ack => W_output_data2_3487_delayed_13_0_3656_inst_req_1); -- 
    sendModule_cp_element_group_335: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_335"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_335 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(335), clk => clk, reset => reset); --
    end block;
    -- CP-element group 336:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 336: predecessors 
    -- CP-element group 336: 	334 
    -- CP-element group 336: successors 
    -- CP-element group 336: marked-successors 
    -- CP-element group 336: 	159 
    -- CP-element group 336: 	334 
    -- CP-element group 336:  members (3) 
      -- CP-element group 336: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_sample_completed_
      -- CP-element group 336: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Sample/ack
      -- CP-element group 336: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Sample/$exit
      -- 
    ack_8014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 336_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3487_delayed_13_0_3656_inst_ack_0, ack => sendModule_CP_6819_elements(336)); -- 
    -- CP-element group 337:  transition  input  bypass  pipeline-parent 
    -- CP-element group 337: predecessors 
    -- CP-element group 337: 	335 
    -- CP-element group 337: successors 
    -- CP-element group 337: 	370 
    -- CP-element group 337:  members (3) 
      -- CP-element group 337: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_update_completed_
      -- CP-element group 337: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Update/ack
      -- CP-element group 337: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3658_Update/$exit
      -- 
    ack_8019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 337_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3487_delayed_13_0_3656_inst_ack_1, ack => sendModule_CP_6819_elements(337)); -- 
    -- CP-element group 338:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 338: predecessors 
    -- CP-element group 338: 	43 
    -- CP-element group 338: marked-predecessors 
    -- CP-element group 338: 	340 
    -- CP-element group 338: successors 
    -- CP-element group 338: 	340 
    -- CP-element group 338:  members (3) 
      -- CP-element group 338: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Sample/rr
      -- CP-element group 338: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Sample/$entry
      -- CP-element group 338: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_sample_start_
      -- 
    rr_8027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(338), ack => EQ_u3_u1_3668_inst_req_0); -- 
    sendModule_cp_element_group_338: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_338"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(340);
      gj_sendModule_cp_element_group_338 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(338), clk => clk, reset => reset); --
    end block;
    -- CP-element group 339:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 339: predecessors 
    -- CP-element group 339: marked-predecessors 
    -- CP-element group 339: 	372 
    -- CP-element group 339: successors 
    -- CP-element group 339: 	341 
    -- CP-element group 339:  members (3) 
      -- CP-element group 339: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Update/cr
      -- CP-element group 339: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Update/$entry
      -- CP-element group 339: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_update_start_
      -- 
    cr_8032_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8032_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(339), ack => EQ_u3_u1_3668_inst_req_1); -- 
    sendModule_cp_element_group_339: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_339"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_339 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(339), clk => clk, reset => reset); --
    end block;
    -- CP-element group 340:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 340: predecessors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: successors 
    -- CP-element group 340: marked-successors 
    -- CP-element group 340: 	338 
    -- CP-element group 340: 	41 
    -- CP-element group 340:  members (3) 
      -- CP-element group 340: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Sample/ra
      -- CP-element group 340: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Sample/$exit
      -- CP-element group 340: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_sample_completed_
      -- 
    ra_8028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 340_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3668_inst_ack_0, ack => sendModule_CP_6819_elements(340)); -- 
    -- CP-element group 341:  transition  input  bypass  pipeline-parent 
    -- CP-element group 341: predecessors 
    -- CP-element group 341: 	339 
    -- CP-element group 341: successors 
    -- CP-element group 341: 	370 
    -- CP-element group 341:  members (3) 
      -- CP-element group 341: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Update/ca
      -- CP-element group 341: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_Update/$exit
      -- CP-element group 341: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3668_update_completed_
      -- 
    ca_8033_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 341_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3668_inst_ack_1, ack => sendModule_CP_6819_elements(341)); -- 
    -- CP-element group 342:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 342: predecessors 
    -- CP-element group 342: 	161 
    -- CP-element group 342: marked-predecessors 
    -- CP-element group 342: 	344 
    -- CP-element group 342: successors 
    -- CP-element group 342: 	344 
    -- CP-element group 342:  members (3) 
      -- CP-element group 342: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_sample_start_
      -- CP-element group 342: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Sample/req
      -- CP-element group 342: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Sample/$entry
      -- 
    req_8041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(342), ack => W_output_data2_3495_delayed_13_0_3670_inst_req_0); -- 
    sendModule_cp_element_group_342: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_342"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(344);
      gj_sendModule_cp_element_group_342 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(342), clk => clk, reset => reset); --
    end block;
    -- CP-element group 343:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 343: predecessors 
    -- CP-element group 343: marked-predecessors 
    -- CP-element group 343: 	372 
    -- CP-element group 343: successors 
    -- CP-element group 343: 	345 
    -- CP-element group 343:  members (3) 
      -- CP-element group 343: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Update/$entry
      -- CP-element group 343: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_update_start_
      -- CP-element group 343: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Update/req
      -- 
    req_8046_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8046_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(343), ack => W_output_data2_3495_delayed_13_0_3670_inst_req_1); -- 
    sendModule_cp_element_group_343: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_343"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_343 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(343), clk => clk, reset => reset); --
    end block;
    -- CP-element group 344:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 344: predecessors 
    -- CP-element group 344: 	342 
    -- CP-element group 344: successors 
    -- CP-element group 344: marked-successors 
    -- CP-element group 344: 	159 
    -- CP-element group 344: 	342 
    -- CP-element group 344:  members (3) 
      -- CP-element group 344: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Sample/ack
      -- CP-element group 344: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_sample_completed_
      -- CP-element group 344: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Sample/$exit
      -- 
    ack_8042_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 344_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3495_delayed_13_0_3670_inst_ack_0, ack => sendModule_CP_6819_elements(344)); -- 
    -- CP-element group 345:  transition  input  bypass  pipeline-parent 
    -- CP-element group 345: predecessors 
    -- CP-element group 345: 	343 
    -- CP-element group 345: successors 
    -- CP-element group 345: 	370 
    -- CP-element group 345:  members (3) 
      -- CP-element group 345: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Update/$exit
      -- CP-element group 345: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_update_completed_
      -- CP-element group 345: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3672_Update/ack
      -- 
    ack_8047_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 345_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3495_delayed_13_0_3670_inst_ack_1, ack => sendModule_CP_6819_elements(345)); -- 
    -- CP-element group 346:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 346: predecessors 
    -- CP-element group 346: 	43 
    -- CP-element group 346: marked-predecessors 
    -- CP-element group 346: 	348 
    -- CP-element group 346: successors 
    -- CP-element group 346: 	348 
    -- CP-element group 346:  members (3) 
      -- CP-element group 346: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Sample/$entry
      -- CP-element group 346: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Sample/rr
      -- CP-element group 346: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_sample_start_
      -- 
    rr_8055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(346), ack => EQ_u3_u1_3682_inst_req_0); -- 
    sendModule_cp_element_group_346: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_346"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(43) & sendModule_CP_6819_elements(348);
      gj_sendModule_cp_element_group_346 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(346), clk => clk, reset => reset); --
    end block;
    -- CP-element group 347:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 347: predecessors 
    -- CP-element group 347: marked-predecessors 
    -- CP-element group 347: 	372 
    -- CP-element group 347: successors 
    -- CP-element group 347: 	349 
    -- CP-element group 347:  members (3) 
      -- CP-element group 347: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Update/cr
      -- CP-element group 347: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Update/$entry
      -- CP-element group 347: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_update_start_
      -- 
    cr_8060_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8060_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(347), ack => EQ_u3_u1_3682_inst_req_1); -- 
    sendModule_cp_element_group_347: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_347"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_347 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(347), clk => clk, reset => reset); --
    end block;
    -- CP-element group 348:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 348: predecessors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: successors 
    -- CP-element group 348: marked-successors 
    -- CP-element group 348: 	346 
    -- CP-element group 348: 	41 
    -- CP-element group 348:  members (3) 
      -- CP-element group 348: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Sample/ra
      -- CP-element group 348: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_sample_completed_
      -- CP-element group 348: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Sample/$exit
      -- 
    ra_8056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 348_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3682_inst_ack_0, ack => sendModule_CP_6819_elements(348)); -- 
    -- CP-element group 349:  transition  input  bypass  pipeline-parent 
    -- CP-element group 349: predecessors 
    -- CP-element group 349: 	347 
    -- CP-element group 349: successors 
    -- CP-element group 349: 	370 
    -- CP-element group 349:  members (3) 
      -- CP-element group 349: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_update_completed_
      -- CP-element group 349: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Update/$exit
      -- CP-element group 349: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/EQ_u3_u1_3682_Update/ca
      -- 
    ca_8061_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 349_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u3_u1_3682_inst_ack_1, ack => sendModule_CP_6819_elements(349)); -- 
    -- CP-element group 350:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 350: predecessors 
    -- CP-element group 350: 	161 
    -- CP-element group 350: marked-predecessors 
    -- CP-element group 350: 	352 
    -- CP-element group 350: successors 
    -- CP-element group 350: 	352 
    -- CP-element group 350:  members (3) 
      -- CP-element group 350: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_sample_start_
      -- CP-element group 350: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Sample/req
      -- CP-element group 350: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Sample/$entry
      -- 
    req_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(350), ack => W_output_data2_3503_delayed_13_0_3684_inst_req_0); -- 
    sendModule_cp_element_group_350: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_350"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(161) & sendModule_CP_6819_elements(352);
      gj_sendModule_cp_element_group_350 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(350), clk => clk, reset => reset); --
    end block;
    -- CP-element group 351:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 351: predecessors 
    -- CP-element group 351: marked-predecessors 
    -- CP-element group 351: 	372 
    -- CP-element group 351: successors 
    -- CP-element group 351: 	353 
    -- CP-element group 351:  members (3) 
      -- CP-element group 351: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_update_start_
      -- CP-element group 351: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Update/$entry
      -- CP-element group 351: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Update/req
      -- 
    req_8074_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8074_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(351), ack => W_output_data2_3503_delayed_13_0_3684_inst_req_1); -- 
    sendModule_cp_element_group_351: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_351"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_351 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(351), clk => clk, reset => reset); --
    end block;
    -- CP-element group 352:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 352: predecessors 
    -- CP-element group 352: 	350 
    -- CP-element group 352: successors 
    -- CP-element group 352: marked-successors 
    -- CP-element group 352: 	159 
    -- CP-element group 352: 	350 
    -- CP-element group 352:  members (3) 
      -- CP-element group 352: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Sample/$exit
      -- CP-element group 352: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_sample_completed_
      -- CP-element group 352: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Sample/ack
      -- 
    ack_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 352_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3503_delayed_13_0_3684_inst_ack_0, ack => sendModule_CP_6819_elements(352)); -- 
    -- CP-element group 353:  transition  input  bypass  pipeline-parent 
    -- CP-element group 353: predecessors 
    -- CP-element group 353: 	351 
    -- CP-element group 353: successors 
    -- CP-element group 353: 	370 
    -- CP-element group 353:  members (3) 
      -- CP-element group 353: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_update_completed_
      -- CP-element group 353: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Update/ack
      -- CP-element group 353: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3686_Update/$exit
      -- 
    ack_8075_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 353_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_output_data2_3503_delayed_13_0_3684_inst_ack_1, ack => sendModule_CP_6819_elements(353)); -- 
    -- CP-element group 354:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 354: predecessors 
    -- CP-element group 354: 	134 
    -- CP-element group 354: marked-predecessors 
    -- CP-element group 354: 	356 
    -- CP-element group 354: successors 
    -- CP-element group 354: 	356 
    -- CP-element group 354:  members (3) 
      -- CP-element group 354: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_sample_start_
      -- CP-element group 354: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Sample/$entry
      -- CP-element group 354: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Sample/req
      -- 
    req_8083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(354), ack => W_fetch_addr1_3507_delayed_8_0_3693_inst_req_0); -- 
    sendModule_cp_element_group_354: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_354"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(134) & sendModule_CP_6819_elements(356);
      gj_sendModule_cp_element_group_354 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(354), clk => clk, reset => reset); --
    end block;
    -- CP-element group 355:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 355: predecessors 
    -- CP-element group 355: marked-predecessors 
    -- CP-element group 355: 	364 
    -- CP-element group 355: successors 
    -- CP-element group 355: 	357 
    -- CP-element group 355:  members (3) 
      -- CP-element group 355: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_update_start_
      -- CP-element group 355: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Update/$entry
      -- CP-element group 355: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Update/req
      -- 
    req_8088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(355), ack => W_fetch_addr1_3507_delayed_8_0_3693_inst_req_1); -- 
    sendModule_cp_element_group_355: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_355"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(364);
      gj_sendModule_cp_element_group_355 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(355), clk => clk, reset => reset); --
    end block;
    -- CP-element group 356:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 356: predecessors 
    -- CP-element group 356: 	354 
    -- CP-element group 356: successors 
    -- CP-element group 356: marked-successors 
    -- CP-element group 356: 	129 
    -- CP-element group 356: 	354 
    -- CP-element group 356:  members (3) 
      -- CP-element group 356: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_sample_completed_
      -- CP-element group 356: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Sample/$exit
      -- CP-element group 356: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Sample/ack
      -- 
    ack_8084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 356_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_0, ack => sendModule_CP_6819_elements(356)); -- 
    -- CP-element group 357:  transition  input  bypass  pipeline-parent 
    -- CP-element group 357: predecessors 
    -- CP-element group 357: 	355 
    -- CP-element group 357: successors 
    -- CP-element group 357: 	362 
    -- CP-element group 357:  members (19) 
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_update_completed_
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Update/$exit
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3695_Update/ack
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_word_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_root_address_calculated
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_address_resized
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_addr_resize/$entry
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_addr_resize/$exit
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_addr_resize/base_resize_req
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_addr_resize/base_resize_ack
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_plus_offset/$entry
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_plus_offset/$exit
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_plus_offset/sum_rename_req
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_base_plus_offset/sum_rename_ack
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_word_addrgen/$entry
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_word_addrgen/$exit
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_word_addrgen/root_register_req
      -- CP-element group 357: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_word_addrgen/root_register_ack
      -- 
    ack_8089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 357_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_1, ack => sendModule_CP_6819_elements(357)); -- 
    -- CP-element group 358:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 358: predecessors 
    -- CP-element group 358: 	165 
    -- CP-element group 358: 	169 
    -- CP-element group 358: 	173 
    -- CP-element group 358: 	177 
    -- CP-element group 358: 	181 
    -- CP-element group 358: 	185 
    -- CP-element group 358: 	189 
    -- CP-element group 358: 	193 
    -- CP-element group 358: 	229 
    -- CP-element group 358: 	233 
    -- CP-element group 358: 	237 
    -- CP-element group 358: 	241 
    -- CP-element group 358: 	245 
    -- CP-element group 358: 	249 
    -- CP-element group 358: 	253 
    -- CP-element group 358: 	257 
    -- CP-element group 358: 	261 
    -- CP-element group 358: 	265 
    -- CP-element group 358: 	269 
    -- CP-element group 358: 	273 
    -- CP-element group 358: 	277 
    -- CP-element group 358: 	281 
    -- CP-element group 358: 	285 
    -- CP-element group 358: 	289 
    -- CP-element group 358: marked-predecessors 
    -- CP-element group 358: 	360 
    -- CP-element group 358: successors 
    -- CP-element group 358: 	360 
    -- CP-element group 358:  members (3) 
      -- CP-element group 358: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_sample_start_
      -- CP-element group 358: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Sample/$entry
      -- CP-element group 358: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Sample/rr
      -- 
    rr_8097_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8097_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(358), ack => CONCAT_u32_u64_3712_inst_req_0); -- 
    sendModule_cp_element_group_358: block -- 
      constant place_capacities: IntegerArray(0 to 24) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1);
      constant place_markings: IntegerArray(0 to 24)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant place_delays: IntegerArray(0 to 24) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_358"; 
      signal preds: BooleanArray(1 to 25); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(165) & sendModule_CP_6819_elements(169) & sendModule_CP_6819_elements(173) & sendModule_CP_6819_elements(177) & sendModule_CP_6819_elements(181) & sendModule_CP_6819_elements(185) & sendModule_CP_6819_elements(189) & sendModule_CP_6819_elements(193) & sendModule_CP_6819_elements(229) & sendModule_CP_6819_elements(233) & sendModule_CP_6819_elements(237) & sendModule_CP_6819_elements(241) & sendModule_CP_6819_elements(245) & sendModule_CP_6819_elements(249) & sendModule_CP_6819_elements(253) & sendModule_CP_6819_elements(257) & sendModule_CP_6819_elements(261) & sendModule_CP_6819_elements(265) & sendModule_CP_6819_elements(269) & sendModule_CP_6819_elements(273) & sendModule_CP_6819_elements(277) & sendModule_CP_6819_elements(281) & sendModule_CP_6819_elements(285) & sendModule_CP_6819_elements(289) & sendModule_CP_6819_elements(360);
      gj_sendModule_cp_element_group_358 : generic_join generic map(name => joinName, number_of_predecessors => 25, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(358), clk => clk, reset => reset); --
    end block;
    -- CP-element group 359:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 359: predecessors 
    -- CP-element group 359: marked-predecessors 
    -- CP-element group 359: 	364 
    -- CP-element group 359: successors 
    -- CP-element group 359: 	361 
    -- CP-element group 359:  members (3) 
      -- CP-element group 359: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_update_start_
      -- CP-element group 359: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Update/$entry
      -- CP-element group 359: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Update/cr
      -- 
    cr_8102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(359), ack => CONCAT_u32_u64_3712_inst_req_1); -- 
    sendModule_cp_element_group_359: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_359"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(364);
      gj_sendModule_cp_element_group_359 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(359), clk => clk, reset => reset); --
    end block;
    -- CP-element group 360:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 360: predecessors 
    -- CP-element group 360: 	358 
    -- CP-element group 360: successors 
    -- CP-element group 360: marked-successors 
    -- CP-element group 360: 	163 
    -- CP-element group 360: 	167 
    -- CP-element group 360: 	171 
    -- CP-element group 360: 	175 
    -- CP-element group 360: 	179 
    -- CP-element group 360: 	183 
    -- CP-element group 360: 	187 
    -- CP-element group 360: 	191 
    -- CP-element group 360: 	227 
    -- CP-element group 360: 	231 
    -- CP-element group 360: 	235 
    -- CP-element group 360: 	239 
    -- CP-element group 360: 	243 
    -- CP-element group 360: 	247 
    -- CP-element group 360: 	251 
    -- CP-element group 360: 	255 
    -- CP-element group 360: 	259 
    -- CP-element group 360: 	263 
    -- CP-element group 360: 	267 
    -- CP-element group 360: 	271 
    -- CP-element group 360: 	275 
    -- CP-element group 360: 	279 
    -- CP-element group 360: 	283 
    -- CP-element group 360: 	287 
    -- CP-element group 360: 	358 
    -- CP-element group 360:  members (3) 
      -- CP-element group 360: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_sample_completed_
      -- CP-element group 360: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Sample/$exit
      -- CP-element group 360: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Sample/ra
      -- 
    ra_8098_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 360_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3712_inst_ack_0, ack => sendModule_CP_6819_elements(360)); -- 
    -- CP-element group 361:  transition  input  bypass  pipeline-parent 
    -- CP-element group 361: predecessors 
    -- CP-element group 361: 	359 
    -- CP-element group 361: successors 
    -- CP-element group 361: 	362 
    -- CP-element group 361:  members (3) 
      -- CP-element group 361: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_update_completed_
      -- CP-element group 361: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Update/$exit
      -- CP-element group 361: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3712_Update/ca
      -- 
    ca_8103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 361_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3712_inst_ack_1, ack => sendModule_CP_6819_elements(361)); -- 
    -- CP-element group 362:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 362: predecessors 
    -- CP-element group 362: 	357 
    -- CP-element group 362: 	361 
    -- CP-element group 362: 	383 
    -- CP-element group 362: 	384 
    -- CP-element group 362: marked-predecessors 
    -- CP-element group 362: 	364 
    -- CP-element group 362: successors 
    -- CP-element group 362: 	364 
    -- CP-element group 362:  members (9) 
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_sample_start_
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/$entry
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/ptr_deref_3697_Split/$entry
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/ptr_deref_3697_Split/$exit
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/ptr_deref_3697_Split/split_req
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/ptr_deref_3697_Split/split_ack
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/$entry
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/word_0/$entry
      -- CP-element group 362: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/word_0/rr
      -- 
    rr_8141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(362), ack => ptr_deref_3697_store_0_req_0); -- 
    sendModule_cp_element_group_362: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_362"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(357) & sendModule_CP_6819_elements(361) & sendModule_CP_6819_elements(383) & sendModule_CP_6819_elements(384) & sendModule_CP_6819_elements(364);
      gj_sendModule_cp_element_group_362 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(362), clk => clk, reset => reset); --
    end block;
    -- CP-element group 363:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 363: predecessors 
    -- CP-element group 363: marked-predecessors 
    -- CP-element group 363: 	365 
    -- CP-element group 363: successors 
    -- CP-element group 363: 	365 
    -- CP-element group 363:  members (5) 
      -- CP-element group 363: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_update_start_
      -- CP-element group 363: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/$entry
      -- CP-element group 363: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/$entry
      -- CP-element group 363: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/word_0/$entry
      -- CP-element group 363: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/word_0/cr
      -- 
    cr_8152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(363), ack => ptr_deref_3697_store_0_req_1); -- 
    sendModule_cp_element_group_363: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_363"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(365);
      gj_sendModule_cp_element_group_363 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(363), clk => clk, reset => reset); --
    end block;
    -- CP-element group 364:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 364: predecessors 
    -- CP-element group 364: 	362 
    -- CP-element group 364: successors 
    -- CP-element group 364: 	385 
    -- CP-element group 364: marked-successors 
    -- CP-element group 364: 	355 
    -- CP-element group 364: 	359 
    -- CP-element group 364: 	362 
    -- CP-element group 364:  members (5) 
      -- CP-element group 364: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_sample_completed_
      -- CP-element group 364: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/$exit
      -- CP-element group 364: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/$exit
      -- CP-element group 364: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/word_0/$exit
      -- CP-element group 364: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Sample/word_access_start/word_0/ra
      -- 
    ra_8142_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 364_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3697_store_0_ack_0, ack => sendModule_CP_6819_elements(364)); -- 
    -- CP-element group 365:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 365: predecessors 
    -- CP-element group 365: 	363 
    -- CP-element group 365: successors 
    -- CP-element group 365: 	386 
    -- CP-element group 365: marked-successors 
    -- CP-element group 365: 	363 
    -- CP-element group 365:  members (5) 
      -- CP-element group 365: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_update_completed_
      -- CP-element group 365: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/$exit
      -- CP-element group 365: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/$exit
      -- CP-element group 365: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/word_0/$exit
      -- CP-element group 365: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_Update/word_access_complete/word_0/ca
      -- 
    ca_8153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 365_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3697_store_0_ack_1, ack => sendModule_CP_6819_elements(365)); -- 
    -- CP-element group 366:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 366: predecessors 
    -- CP-element group 366: 	141 
    -- CP-element group 366: marked-predecessors 
    -- CP-element group 366: 	368 
    -- CP-element group 366: successors 
    -- CP-element group 366: 	368 
    -- CP-element group 366:  members (3) 
      -- CP-element group 366: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_sample_start_
      -- CP-element group 366: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Sample/$entry
      -- CP-element group 366: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Sample/req
      -- 
    req_8161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(366), ack => W_fetch_addr2_3525_delayed_8_0_3714_inst_req_0); -- 
    sendModule_cp_element_group_366: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_366"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(141) & sendModule_CP_6819_elements(368);
      gj_sendModule_cp_element_group_366 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(366), clk => clk, reset => reset); --
    end block;
    -- CP-element group 367:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 367: predecessors 
    -- CP-element group 367: marked-predecessors 
    -- CP-element group 367: 	376 
    -- CP-element group 367: successors 
    -- CP-element group 367: 	369 
    -- CP-element group 367:  members (3) 
      -- CP-element group 367: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_update_start_
      -- CP-element group 367: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Update/$entry
      -- CP-element group 367: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Update/req
      -- 
    req_8166_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8166_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(367), ack => W_fetch_addr2_3525_delayed_8_0_3714_inst_req_1); -- 
    sendModule_cp_element_group_367: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_367"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(376);
      gj_sendModule_cp_element_group_367 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(367), clk => clk, reset => reset); --
    end block;
    -- CP-element group 368:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 368: predecessors 
    -- CP-element group 368: 	366 
    -- CP-element group 368: successors 
    -- CP-element group 368: marked-successors 
    -- CP-element group 368: 	136 
    -- CP-element group 368: 	366 
    -- CP-element group 368:  members (3) 
      -- CP-element group 368: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_sample_completed_
      -- CP-element group 368: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Sample/$exit
      -- CP-element group 368: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Sample/ack
      -- 
    ack_8162_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 368_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_0, ack => sendModule_CP_6819_elements(368)); -- 
    -- CP-element group 369:  transition  input  bypass  pipeline-parent 
    -- CP-element group 369: predecessors 
    -- CP-element group 369: 	367 
    -- CP-element group 369: successors 
    -- CP-element group 369: 	374 
    -- CP-element group 369:  members (19) 
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_update_completed_
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Update/$exit
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/assign_stmt_3716_Update/ack
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_word_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_root_address_calculated
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_address_resized
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_addr_resize/$entry
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_addr_resize/$exit
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_addr_resize/base_resize_req
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_addr_resize/base_resize_ack
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_plus_offset/$entry
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_plus_offset/$exit
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_plus_offset/sum_rename_req
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_base_plus_offset/sum_rename_ack
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_word_addrgen/$entry
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_word_addrgen/$exit
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_word_addrgen/root_register_req
      -- CP-element group 369: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_word_addrgen/root_register_ack
      -- 
    ack_8167_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 369_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_1, ack => sendModule_CP_6819_elements(369)); -- 
    -- CP-element group 370:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 370: predecessors 
    -- CP-element group 370: 	197 
    -- CP-element group 370: 	201 
    -- CP-element group 370: 	205 
    -- CP-element group 370: 	209 
    -- CP-element group 370: 	213 
    -- CP-element group 370: 	217 
    -- CP-element group 370: 	221 
    -- CP-element group 370: 	225 
    -- CP-element group 370: 	293 
    -- CP-element group 370: 	297 
    -- CP-element group 370: 	301 
    -- CP-element group 370: 	305 
    -- CP-element group 370: 	309 
    -- CP-element group 370: 	313 
    -- CP-element group 370: 	317 
    -- CP-element group 370: 	321 
    -- CP-element group 370: 	325 
    -- CP-element group 370: 	329 
    -- CP-element group 370: 	333 
    -- CP-element group 370: 	337 
    -- CP-element group 370: 	341 
    -- CP-element group 370: 	345 
    -- CP-element group 370: 	349 
    -- CP-element group 370: 	353 
    -- CP-element group 370: marked-predecessors 
    -- CP-element group 370: 	372 
    -- CP-element group 370: successors 
    -- CP-element group 370: 	372 
    -- CP-element group 370:  members (3) 
      -- CP-element group 370: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_sample_start_
      -- CP-element group 370: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Sample/$entry
      -- CP-element group 370: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Sample/rr
      -- 
    rr_8175_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8175_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(370), ack => CONCAT_u32_u64_3733_inst_req_0); -- 
    sendModule_cp_element_group_370: block -- 
      constant place_capacities: IntegerArray(0 to 24) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1,19 => 1,20 => 1,21 => 1,22 => 1,23 => 1,24 => 1);
      constant place_markings: IntegerArray(0 to 24)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant place_delays: IntegerArray(0 to 24) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0,19 => 0,20 => 0,21 => 0,22 => 0,23 => 0,24 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_370"; 
      signal preds: BooleanArray(1 to 25); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(197) & sendModule_CP_6819_elements(201) & sendModule_CP_6819_elements(205) & sendModule_CP_6819_elements(209) & sendModule_CP_6819_elements(213) & sendModule_CP_6819_elements(217) & sendModule_CP_6819_elements(221) & sendModule_CP_6819_elements(225) & sendModule_CP_6819_elements(293) & sendModule_CP_6819_elements(297) & sendModule_CP_6819_elements(301) & sendModule_CP_6819_elements(305) & sendModule_CP_6819_elements(309) & sendModule_CP_6819_elements(313) & sendModule_CP_6819_elements(317) & sendModule_CP_6819_elements(321) & sendModule_CP_6819_elements(325) & sendModule_CP_6819_elements(329) & sendModule_CP_6819_elements(333) & sendModule_CP_6819_elements(337) & sendModule_CP_6819_elements(341) & sendModule_CP_6819_elements(345) & sendModule_CP_6819_elements(349) & sendModule_CP_6819_elements(353) & sendModule_CP_6819_elements(372);
      gj_sendModule_cp_element_group_370 : generic_join generic map(name => joinName, number_of_predecessors => 25, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(370), clk => clk, reset => reset); --
    end block;
    -- CP-element group 371:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 371: predecessors 
    -- CP-element group 371: marked-predecessors 
    -- CP-element group 371: 	376 
    -- CP-element group 371: successors 
    -- CP-element group 371: 	373 
    -- CP-element group 371:  members (3) 
      -- CP-element group 371: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_update_start_
      -- CP-element group 371: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Update/$entry
      -- CP-element group 371: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Update/cr
      -- 
    cr_8180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(371), ack => CONCAT_u32_u64_3733_inst_req_1); -- 
    sendModule_cp_element_group_371: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_371"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(376);
      gj_sendModule_cp_element_group_371 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(371), clk => clk, reset => reset); --
    end block;
    -- CP-element group 372:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 372: predecessors 
    -- CP-element group 372: 	370 
    -- CP-element group 372: successors 
    -- CP-element group 372: marked-successors 
    -- CP-element group 372: 	195 
    -- CP-element group 372: 	199 
    -- CP-element group 372: 	203 
    -- CP-element group 372: 	207 
    -- CP-element group 372: 	211 
    -- CP-element group 372: 	215 
    -- CP-element group 372: 	219 
    -- CP-element group 372: 	223 
    -- CP-element group 372: 	291 
    -- CP-element group 372: 	295 
    -- CP-element group 372: 	299 
    -- CP-element group 372: 	303 
    -- CP-element group 372: 	307 
    -- CP-element group 372: 	311 
    -- CP-element group 372: 	315 
    -- CP-element group 372: 	319 
    -- CP-element group 372: 	323 
    -- CP-element group 372: 	327 
    -- CP-element group 372: 	331 
    -- CP-element group 372: 	335 
    -- CP-element group 372: 	339 
    -- CP-element group 372: 	343 
    -- CP-element group 372: 	347 
    -- CP-element group 372: 	351 
    -- CP-element group 372: 	370 
    -- CP-element group 372:  members (3) 
      -- CP-element group 372: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_sample_completed_
      -- CP-element group 372: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Sample/$exit
      -- CP-element group 372: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Sample/ra
      -- 
    ra_8176_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 372_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3733_inst_ack_0, ack => sendModule_CP_6819_elements(372)); -- 
    -- CP-element group 373:  transition  input  bypass  pipeline-parent 
    -- CP-element group 373: predecessors 
    -- CP-element group 373: 	371 
    -- CP-element group 373: successors 
    -- CP-element group 373: 	374 
    -- CP-element group 373:  members (3) 
      -- CP-element group 373: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_update_completed_
      -- CP-element group 373: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Update/$exit
      -- CP-element group 373: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/CONCAT_u32_u64_3733_Update/ca
      -- 
    ca_8181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 373_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u32_u64_3733_inst_ack_1, ack => sendModule_CP_6819_elements(373)); -- 
    -- CP-element group 374:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 374: predecessors 
    -- CP-element group 374: 	369 
    -- CP-element group 374: 	373 
    -- CP-element group 374: 	385 
    -- CP-element group 374: marked-predecessors 
    -- CP-element group 374: 	376 
    -- CP-element group 374: successors 
    -- CP-element group 374: 	376 
    -- CP-element group 374:  members (9) 
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_sample_start_
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/$entry
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/ptr_deref_3718_Split/$entry
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/ptr_deref_3718_Split/$exit
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/ptr_deref_3718_Split/split_req
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/ptr_deref_3718_Split/split_ack
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/$entry
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/word_0/$entry
      -- CP-element group 374: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/word_0/rr
      -- 
    rr_8219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(374), ack => ptr_deref_3718_store_0_req_0); -- 
    sendModule_cp_element_group_374: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_374"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(369) & sendModule_CP_6819_elements(373) & sendModule_CP_6819_elements(385) & sendModule_CP_6819_elements(376);
      gj_sendModule_cp_element_group_374 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(374), clk => clk, reset => reset); --
    end block;
    -- CP-element group 375:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 375: predecessors 
    -- CP-element group 375: marked-predecessors 
    -- CP-element group 375: 	377 
    -- CP-element group 375: successors 
    -- CP-element group 375: 	377 
    -- CP-element group 375:  members (5) 
      -- CP-element group 375: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_update_start_
      -- CP-element group 375: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/$entry
      -- CP-element group 375: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/$entry
      -- CP-element group 375: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/word_0/$entry
      -- CP-element group 375: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/word_0/cr
      -- 
    cr_8230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(375), ack => ptr_deref_3718_store_0_req_1); -- 
    sendModule_cp_element_group_375: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_375"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(377);
      gj_sendModule_cp_element_group_375 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(375), clk => clk, reset => reset); --
    end block;
    -- CP-element group 376:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 376: predecessors 
    -- CP-element group 376: 	374 
    -- CP-element group 376: successors 
    -- CP-element group 376: 	386 
    -- CP-element group 376: marked-successors 
    -- CP-element group 376: 	142 
    -- CP-element group 376: 	146 
    -- CP-element group 376: 	367 
    -- CP-element group 376: 	371 
    -- CP-element group 376: 	374 
    -- CP-element group 376:  members (6) 
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_sample_completed_
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/$exit
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/$exit
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/word_0/$exit
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Sample/word_access_start/word_0/ra
      -- CP-element group 376: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ring_reenable_memory_space_0
      -- 
    ra_8220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 376_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3718_store_0_ack_0, ack => sendModule_CP_6819_elements(376)); -- 
    -- CP-element group 377:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 377: predecessors 
    -- CP-element group 377: 	375 
    -- CP-element group 377: successors 
    -- CP-element group 377: 	386 
    -- CP-element group 377: marked-successors 
    -- CP-element group 377: 	375 
    -- CP-element group 377:  members (5) 
      -- CP-element group 377: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_update_completed_
      -- CP-element group 377: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/$exit
      -- CP-element group 377: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/$exit
      -- CP-element group 377: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/word_0/$exit
      -- CP-element group 377: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3718_Update/word_access_complete/word_0/ca
      -- 
    ca_8231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 377_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3718_store_0_ack_1, ack => sendModule_CP_6819_elements(377)); -- 
    -- CP-element group 378:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 378: predecessors 
    -- CP-element group 378: 	15 
    -- CP-element group 378: marked-predecessors 
    -- CP-element group 378: 	380 
    -- CP-element group 378: successors 
    -- CP-element group 378: 	380 
    -- CP-element group 378:  members (3) 
      -- CP-element group 378: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_sample_start_
      -- CP-element group 378: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Sample/$entry
      -- CP-element group 378: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Sample/rr
      -- 
    rr_8239_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8239_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(378), ack => SUB_u16_u16_3738_inst_req_0); -- 
    sendModule_cp_element_group_378: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_378"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(15) & sendModule_CP_6819_elements(380);
      gj_sendModule_cp_element_group_378 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(378), clk => clk, reset => reset); --
    end block;
    -- CP-element group 379:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 379: predecessors 
    -- CP-element group 379: marked-predecessors 
    -- CP-element group 379: 	381 
    -- CP-element group 379: successors 
    -- CP-element group 379: 	381 
    -- CP-element group 379:  members (3) 
      -- CP-element group 379: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_update_start_
      -- CP-element group 379: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Update/$entry
      -- CP-element group 379: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Update/cr
      -- 
    cr_8244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(379), ack => SUB_u16_u16_3738_inst_req_1); -- 
    sendModule_cp_element_group_379: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_379"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= sendModule_CP_6819_elements(381);
      gj_sendModule_cp_element_group_379 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(379), clk => clk, reset => reset); --
    end block;
    -- CP-element group 380:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 380: predecessors 
    -- CP-element group 380: 	378 
    -- CP-element group 380: successors 
    -- CP-element group 380: marked-successors 
    -- CP-element group 380: 	378 
    -- CP-element group 380:  members (3) 
      -- CP-element group 380: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_sample_completed_
      -- CP-element group 380: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Sample/$exit
      -- CP-element group 380: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Sample/ra
      -- 
    ra_8240_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 380_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3738_inst_ack_0, ack => sendModule_CP_6819_elements(380)); -- 
    -- CP-element group 381:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 381: predecessors 
    -- CP-element group 381: 	379 
    -- CP-element group 381: successors 
    -- CP-element group 381: 	16 
    -- CP-element group 381: marked-successors 
    -- CP-element group 381: 	379 
    -- CP-element group 381:  members (3) 
      -- CP-element group 381: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_update_completed_
      -- CP-element group 381: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Update/$exit
      -- CP-element group 381: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/SUB_u16_u16_3738_Update/ca
      -- 
    ca_8245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 381_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u16_u16_3738_inst_ack_1, ack => sendModule_CP_6819_elements(381)); -- 
    -- CP-element group 382:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 382: predecessors 
    -- CP-element group 382: 	15 
    -- CP-element group 382: successors 
    -- CP-element group 382: 	16 
    -- CP-element group 382:  members (1) 
      -- CP-element group 382: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group sendModule_CP_6819_elements(382) is a control-delay.
    cp_element_382_delay: control_delay_element  generic map(name => " 382_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(15), ack => sendModule_CP_6819_elements(382), clk => clk, reset =>reset);
    -- CP-element group 383:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 383: predecessors 
    -- CP-element group 383: 	144 
    -- CP-element group 383: successors 
    -- CP-element group 383: 	362 
    -- CP-element group 383:  members (1) 
      -- CP-element group 383: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3380_ptr_deref_3697_delay
      -- 
    -- Element group sendModule_CP_6819_elements(383) is a control-delay.
    cp_element_383_delay: control_delay_element  generic map(name => " 383_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(144), ack => sendModule_CP_6819_elements(383), clk => clk, reset =>reset);
    -- CP-element group 384:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 384: predecessors 
    -- CP-element group 384: 	148 
    -- CP-element group 384: successors 
    -- CP-element group 384: 	362 
    -- CP-element group 384:  members (1) 
      -- CP-element group 384: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3384_ptr_deref_3697_delay
      -- 
    -- Element group sendModule_CP_6819_elements(384) is a control-delay.
    cp_element_384_delay: control_delay_element  generic map(name => " 384_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(148), ack => sendModule_CP_6819_elements(384), clk => clk, reset =>reset);
    -- CP-element group 385:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 385: predecessors 
    -- CP-element group 385: 	364 
    -- CP-element group 385: successors 
    -- CP-element group 385: 	374 
    -- CP-element group 385:  members (1) 
      -- CP-element group 385: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/ptr_deref_3697_ptr_deref_3718_delay
      -- 
    -- Element group sendModule_CP_6819_elements(385) is a control-delay.
    cp_element_385_delay: control_delay_element  generic map(name => " 385_delay", delay_value => 1)  port map(req => sendModule_CP_6819_elements(364), ack => sendModule_CP_6819_elements(385), clk => clk, reset =>reset);
    -- CP-element group 386:  join  transition  bypass  pipeline-parent 
    -- CP-element group 386: predecessors 
    -- CP-element group 386: 	123 
    -- CP-element group 386: 	127 
    -- CP-element group 386: 	131 
    -- CP-element group 386: 	138 
    -- CP-element group 386: 	365 
    -- CP-element group 386: 	376 
    -- CP-element group 386: 	377 
    -- CP-element group 386: 	18 
    -- CP-element group 386: successors 
    -- CP-element group 386: 	12 
    -- CP-element group 386:  members (1) 
      -- CP-element group 386: 	 branch_block_stmt_3226/do_while_stmt_3242/do_while_stmt_3242_loop_body/$exit
      -- 
    sendModule_cp_element_group_386: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 31) := "sendModule_cp_element_group_386"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= sendModule_CP_6819_elements(123) & sendModule_CP_6819_elements(127) & sendModule_CP_6819_elements(131) & sendModule_CP_6819_elements(138) & sendModule_CP_6819_elements(365) & sendModule_CP_6819_elements(376) & sendModule_CP_6819_elements(377) & sendModule_CP_6819_elements(18);
      gj_sendModule_cp_element_group_386 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendModule_CP_6819_elements(386), clk => clk, reset => reset); --
    end block;
    -- CP-element group 387:  transition  input  bypass  pipeline-parent 
    -- CP-element group 387: predecessors 
    -- CP-element group 387: 	11 
    -- CP-element group 387: successors 
    -- CP-element group 387:  members (2) 
      -- CP-element group 387: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_exit/$exit
      -- CP-element group 387: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_exit/ack
      -- 
    ack_8254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 387_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3242_branch_ack_0, ack => sendModule_CP_6819_elements(387)); -- 
    -- CP-element group 388:  transition  input  bypass  pipeline-parent 
    -- CP-element group 388: predecessors 
    -- CP-element group 388: 	11 
    -- CP-element group 388: successors 
    -- CP-element group 388:  members (2) 
      -- CP-element group 388: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_taken/$exit
      -- CP-element group 388: 	 branch_block_stmt_3226/do_while_stmt_3242/loop_taken/ack
      -- 
    ack_8258_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 388_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3242_branch_ack_1, ack => sendModule_CP_6819_elements(388)); -- 
    -- CP-element group 389:  transition  bypass  pipeline-parent 
    -- CP-element group 389: predecessors 
    -- CP-element group 389: 	9 
    -- CP-element group 389: successors 
    -- CP-element group 389: 	1 
    -- CP-element group 389:  members (1) 
      -- CP-element group 389: 	 branch_block_stmt_3226/do_while_stmt_3242/$exit
      -- 
    sendModule_CP_6819_elements(389) <= sendModule_CP_6819_elements(9);
    -- CP-element group 390:  transition  input  output  bypass 
    -- CP-element group 390: predecessors 
    -- CP-element group 390: 	1 
    -- CP-element group 390: successors 
    -- CP-element group 390: 	391 
    -- CP-element group 390:  members (6) 
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_sample_completed_
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_update_start_
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Sample/$exit
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Sample/ack
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Update/$entry
      -- CP-element group 390: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Update/req
      -- 
    ack_8271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 390_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3750_inst_ack_0, ack => sendModule_CP_6819_elements(390)); -- 
    req_8275_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8275_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendModule_CP_6819_elements(390), ack => WPIPE_input_done_pipe_3750_inst_req_1); -- 
    -- CP-element group 391:  transition  place  input  bypass 
    -- CP-element group 391: predecessors 
    -- CP-element group 391: 	390 
    -- CP-element group 391: successors 
    -- CP-element group 391:  members (8) 
      -- CP-element group 391: 	 $exit
      -- CP-element group 391: 	 branch_block_stmt_3226/$exit
      -- CP-element group 391: 	 branch_block_stmt_3226/branch_block_stmt_3226__exit__
      -- CP-element group 391: 	 branch_block_stmt_3226/assign_stmt_3752__exit__
      -- CP-element group 391: 	 branch_block_stmt_3226/assign_stmt_3752/$exit
      -- CP-element group 391: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_update_completed_
      -- CP-element group 391: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Update/$exit
      -- CP-element group 391: 	 branch_block_stmt_3226/assign_stmt_3752/WPIPE_input_done_pipe_3750_Update/ack
      -- 
    ack_8276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 391_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_input_done_pipe_3750_inst_ack_1, ack => sendModule_CP_6819_elements(391)); -- 
    sendModule_do_while_stmt_3242_terminator_8259: loop_terminator -- 
      generic map (name => " sendModule_do_while_stmt_3242_terminator_8259", max_iterations_in_flight =>15) 
      port map(loop_body_exit => sendModule_CP_6819_elements(12),loop_continue => sendModule_CP_6819_elements(388),loop_terminate => sendModule_CP_6819_elements(387),loop_back => sendModule_CP_6819_elements(10),loop_exit => sendModule_CP_6819_elements(9),clk => clk, reset => reset); -- 
    phi_stmt_3244_phi_seq_6941_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_6819_elements(29);
      sendModule_CP_6819_elements(32)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_6819_elements(32);
      sendModule_CP_6819_elements(33)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_6819_elements(34);
      sendModule_CP_6819_elements(30) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_6819_elements(27);
      sendModule_CP_6819_elements(36)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_6819_elements(38);
      sendModule_CP_6819_elements(37)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_6819_elements(39);
      sendModule_CP_6819_elements(28) <= phi_mux_reqs(1);
      phi_stmt_3244_phi_seq_6941 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3244_phi_seq_6941") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_6819_elements(23), 
          phi_sample_ack => sendModule_CP_6819_elements(24), 
          phi_update_req => sendModule_CP_6819_elements(25), 
          phi_update_ack => sendModule_CP_6819_elements(26), 
          phi_mux_ack => sendModule_CP_6819_elements(31), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3249_phi_seq_6995_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_6819_elements(46);
      sendModule_CP_6819_elements(49)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_6819_elements(53);
      sendModule_CP_6819_elements(50)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_6819_elements(54);
      sendModule_CP_6819_elements(47) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_6819_elements(44);
      sendModule_CP_6819_elements(55)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_6819_elements(57);
      sendModule_CP_6819_elements(56)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_6819_elements(58);
      sendModule_CP_6819_elements(45) <= phi_mux_reqs(1);
      phi_stmt_3249_phi_seq_6995 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3249_phi_seq_6995") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_6819_elements(17), 
          phi_sample_ack => sendModule_CP_6819_elements(42), 
          phi_update_req => sendModule_CP_6819_elements(19), 
          phi_update_ack => sendModule_CP_6819_elements(43), 
          phi_mux_ack => sendModule_CP_6819_elements(48), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3254_phi_seq_7039_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_6819_elements(67);
      sendModule_CP_6819_elements(70)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_6819_elements(70);
      sendModule_CP_6819_elements(71)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_6819_elements(72);
      sendModule_CP_6819_elements(68) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_6819_elements(65);
      sendModule_CP_6819_elements(74)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_6819_elements(76);
      sendModule_CP_6819_elements(75)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_6819_elements(77);
      sendModule_CP_6819_elements(66) <= phi_mux_reqs(1);
      phi_stmt_3254_phi_seq_7039 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3254_phi_seq_7039") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_6819_elements(61), 
          phi_sample_ack => sendModule_CP_6819_elements(62), 
          phi_update_req => sendModule_CP_6819_elements(63), 
          phi_update_ack => sendModule_CP_6819_elements(64), 
          phi_mux_ack => sendModule_CP_6819_elements(69), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3259_phi_seq_7083_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_6819_elements(86);
      sendModule_CP_6819_elements(89)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_6819_elements(89);
      sendModule_CP_6819_elements(90)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_6819_elements(91);
      sendModule_CP_6819_elements(87) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_6819_elements(84);
      sendModule_CP_6819_elements(93)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_6819_elements(95);
      sendModule_CP_6819_elements(94)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_6819_elements(96);
      sendModule_CP_6819_elements(85) <= phi_mux_reqs(1);
      phi_stmt_3259_phi_seq_7083 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3259_phi_seq_7083") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_6819_elements(80), 
          phi_sample_ack => sendModule_CP_6819_elements(81), 
          phi_update_req => sendModule_CP_6819_elements(82), 
          phi_update_ack => sendModule_CP_6819_elements(83), 
          phi_mux_ack => sendModule_CP_6819_elements(88), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3264_phi_seq_7127_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= sendModule_CP_6819_elements(105);
      sendModule_CP_6819_elements(108)<= src_sample_reqs(0);
      src_sample_acks(0)  <= sendModule_CP_6819_elements(108);
      sendModule_CP_6819_elements(109)<= src_update_reqs(0);
      src_update_acks(0)  <= sendModule_CP_6819_elements(110);
      sendModule_CP_6819_elements(106) <= phi_mux_reqs(0);
      triggers(1)  <= sendModule_CP_6819_elements(103);
      sendModule_CP_6819_elements(112)<= src_sample_reqs(1);
      src_sample_acks(1)  <= sendModule_CP_6819_elements(114);
      sendModule_CP_6819_elements(113)<= src_update_reqs(1);
      src_update_acks(1)  <= sendModule_CP_6819_elements(115);
      sendModule_CP_6819_elements(104) <= phi_mux_reqs(1);
      phi_stmt_3264_phi_seq_7127 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3264_phi_seq_7127") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => sendModule_CP_6819_elements(99), 
          phi_sample_ack => sendModule_CP_6819_elements(100), 
          phi_update_req => sendModule_CP_6819_elements(101), 
          phi_update_ack => sendModule_CP_6819_elements(102), 
          phi_mux_ack => sendModule_CP_6819_elements(107), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_6893_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= sendModule_CP_6819_elements(13);
        preds(1)  <= sendModule_CP_6819_elements(14);
        entry_tmerge_6893 : transition_merge -- 
          generic map(name => " entry_tmerge_6893")
          port map (preds => preds, symbol_out => sendModule_CP_6819_elements(15));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u16_u16_3292_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3301_wire : std_logic_vector(15 downto 0);
    signal ADD_u16_u16_3310_wire : std_logic_vector(15 downto 0);
    signal ADD_u32_u32_3339_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3349_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_3353_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3704_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3711_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3725_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_3732_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u32_u64_3712_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_3733_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u8_u16_3700_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3703_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3707_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3710_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3721_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3724_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3728_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_3731_wire : std_logic_vector(15 downto 0);
    signal EQ_u3_u1_3382_3382_delayed_14_0_3473 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3390_3390_delayed_14_0_3487 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3398_3398_delayed_14_0_3501 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3406_3406_delayed_14_0_3515 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3414_3414_delayed_14_0_3529 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3422_3422_delayed_14_0_3543 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3430_3430_delayed_14_0_3557 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3438_3438_delayed_14_0_3571 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3446_3446_delayed_14_0_3585 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3454_3454_delayed_14_0_3599 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3462_3462_delayed_14_0_3613 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3470_3470_delayed_14_0_3627 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3478_3478_delayed_14_0_3641 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3486_3486_delayed_14_0_3655 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3494_3494_delayed_14_0_3669 : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_3502_3502_delayed_14_0_3683 : std_logic_vector(0 downto 0);
    signal LSHR_u32_u32_3363_wire : std_logic_vector(31 downto 0);
    signal LSHR_u32_u32_3373_wire : std_logic_vector(31 downto 0);
    signal MUL_u16_u16_3239_wire : std_logic_vector(15 downto 0);
    signal MUX_3303_wire : std_logic_vector(15 downto 0);
    signal MUX_3341_wire : std_logic_vector(31 downto 0);
    signal MUX_3355_wire : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_3745_wire : std_logic_vector(0 downto 0);
    signal SUB_u16_u16_3199_3199_delayed_1_0_3279 : std_logic_vector(15 downto 0);
    signal SUB_u16_u16_3547_3547_delayed_1_0_3739 : std_logic_vector(15 downto 0);
    signal UGE_u16_u1_3284_wire : std_logic_vector(0 downto 0);
    signal ULT_u16_u1_3743_wire : std_logic_vector(0 downto 0);
    signal address1_3244 : std_logic_vector(31 downto 0);
    signal address2_3249 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3365_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3365_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3365_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3365_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3365_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3365_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3375_root_address : std_logic_vector(13 downto 0);
    signal cb_3232 : std_logic_vector(15 downto 0);
    signal chl_3254 : std_logic_vector(15 downto 0);
    signal chl_change_3286 : std_logic_vector(0 downto 0);
    signal chl_out_3235 : std_logic_vector(15 downto 0);
    signal col_3259 : std_logic_vector(15 downto 0);
    signal continue_flag_3747 : std_logic_vector(0 downto 0);
    signal fetch_addr1_3367 : std_logic_vector(31 downto 0);
    signal fetch_addr1_3507_delayed_8_0_3695 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3377 : std_logic_vector(31 downto 0);
    signal fetch_addr2_3525_delayed_8_0_3716 : std_logic_vector(31 downto 0);
    signal fetch_val1_3381 : std_logic_vector(63 downto 0);
    signal fetch_val2_3385 : std_logic_vector(63 downto 0);
    signal konst_3277_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3289_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3291_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3297_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3300_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3309_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3362_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3372_wire_constant : std_logic_vector(31 downto 0);
    signal konst_3471_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3485_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3499_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3513_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3527_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3541_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3555_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3569_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3583_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3597_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3611_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3625_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3639_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3653_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3667_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3681_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3737_wire_constant : std_logic_vector(15 downto 0);
    signal konst_3751_wire_constant : std_logic_vector(7 downto 0);
    signal location1_3464 : std_logic_vector(2 downto 0);
    signal location2_3468 : std_logic_vector(2 downto 0);
    signal n_address1_3343 : std_logic_vector(31 downto 0);
    signal n_address1_3343_3248_buffered : std_logic_vector(31 downto 0);
    signal n_address2_3357 : std_logic_vector(31 downto 0);
    signal n_address2_3357_3253_buffered : std_logic_vector(31 downto 0);
    signal n_chl_3313 : std_logic_vector(15 downto 0);
    signal n_chl_3313_3258_buffered : std_logic_vector(15 downto 0);
    signal n_col_3294 : std_logic_vector(15 downto 0);
    signal n_col_3294_3263_buffered : std_logic_vector(15 downto 0);
    signal n_row_3305 : std_logic_vector(15 downto 0);
    signal n_row_3305_3268_buffered : std_logic_vector(15 downto 0);
    signal output_data1_3383_delayed_13_0_3476 : std_logic_vector(7 downto 0);
    signal output_data1_3391_delayed_13_0_3490 : std_logic_vector(7 downto 0);
    signal output_data1_3392 : std_logic_vector(7 downto 0);
    signal output_data1_3399_delayed_13_0_3504 : std_logic_vector(7 downto 0);
    signal output_data1_3407_delayed_13_0_3518 : std_logic_vector(7 downto 0);
    signal output_data1_3415_delayed_13_0_3532 : std_logic_vector(7 downto 0);
    signal output_data1_3423_delayed_13_0_3546 : std_logic_vector(7 downto 0);
    signal output_data1_3431_delayed_13_0_3560 : std_logic_vector(7 downto 0);
    signal output_data1_3439_delayed_13_0_3574 : std_logic_vector(7 downto 0);
    signal output_data2_3396 : std_logic_vector(7 downto 0);
    signal output_data2_3447_delayed_13_0_3588 : std_logic_vector(7 downto 0);
    signal output_data2_3455_delayed_13_0_3602 : std_logic_vector(7 downto 0);
    signal output_data2_3463_delayed_13_0_3616 : std_logic_vector(7 downto 0);
    signal output_data2_3471_delayed_13_0_3630 : std_logic_vector(7 downto 0);
    signal output_data2_3479_delayed_13_0_3644 : std_logic_vector(7 downto 0);
    signal output_data2_3487_delayed_13_0_3658 : std_logic_vector(7 downto 0);
    signal output_data2_3495_delayed_13_0_3672 : std_logic_vector(7 downto 0);
    signal output_data2_3503_delayed_13_0_3686 : std_logic_vector(7 downto 0);
    signal output_data_read_3388 : std_logic_vector(15 downto 0);
    signal ptr_deref_3380_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3380_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3380_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3380_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3380_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3384_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3384_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3384_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3384_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3384_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3697_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3697_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3697_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3697_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3697_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3697_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3718_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3718_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3718_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3718_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3718_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3718_word_offset_0 : std_logic_vector(13 downto 0);
    signal rb_3229 : std_logic_vector(15 downto 0);
    signal row_3264 : std_logic_vector(15 downto 0);
    signal row_change_3274 : std_logic_vector(0 downto 0);
    signal row_size_3241 : std_logic_vector(31 downto 0);
    signal tmp1_3322 : std_logic_vector(31 downto 0);
    signal tmp2_3331 : std_logic_vector(31 downto 0);
    signal type_cast_3233_3233_delayed_1_0_3317 : std_logic_vector(31 downto 0);
    signal type_cast_3239_3239_delayed_1_0_3326 : std_logic_vector(31 downto 0);
    signal type_cast_3247_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3252_wire : std_logic_vector(31 downto 0);
    signal type_cast_3257_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3262_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3267_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3335_wire : std_logic_vector(31 downto 0);
    signal type_cast_3347_wire : std_logic_vector(31 downto 0);
    signal type_cast_3364_resized : std_logic_vector(13 downto 0);
    signal type_cast_3364_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3364_wire : std_logic_vector(63 downto 0);
    signal type_cast_3374_resized : std_logic_vector(13 downto 0);
    signal type_cast_3374_scaled : std_logic_vector(13 downto 0);
    signal type_cast_3374_wire : std_logic_vector(63 downto 0);
    signal w11_3400 : std_logic_vector(7 downto 0);
    signal w12_3404 : std_logic_vector(7 downto 0);
    signal w13_3408 : std_logic_vector(7 downto 0);
    signal w14_3412 : std_logic_vector(7 downto 0);
    signal w15_3416 : std_logic_vector(7 downto 0);
    signal w16_3420 : std_logic_vector(7 downto 0);
    signal w17_3424 : std_logic_vector(7 downto 0);
    signal w18_3428 : std_logic_vector(7 downto 0);
    signal w21_3432 : std_logic_vector(7 downto 0);
    signal w22_3436 : std_logic_vector(7 downto 0);
    signal w23_3440 : std_logic_vector(7 downto 0);
    signal w24_3444 : std_logic_vector(7 downto 0);
    signal w25_3448 : std_logic_vector(7 downto 0);
    signal w26_3452 : std_logic_vector(7 downto 0);
    signal w27_3456 : std_logic_vector(7 downto 0);
    signal w28_3460 : std_logic_vector(7 downto 0);
    signal wb11_3482 : std_logic_vector(7 downto 0);
    signal wb12_3496 : std_logic_vector(7 downto 0);
    signal wb13_3510 : std_logic_vector(7 downto 0);
    signal wb14_3524 : std_logic_vector(7 downto 0);
    signal wb15_3538 : std_logic_vector(7 downto 0);
    signal wb16_3552 : std_logic_vector(7 downto 0);
    signal wb17_3566 : std_logic_vector(7 downto 0);
    signal wb18_3580 : std_logic_vector(7 downto 0);
    signal wb21_3594 : std_logic_vector(7 downto 0);
    signal wb22_3608 : std_logic_vector(7 downto 0);
    signal wb23_3622 : std_logic_vector(7 downto 0);
    signal wb24_3636 : std_logic_vector(7 downto 0);
    signal wb25_3650 : std_logic_vector(7 downto 0);
    signal wb26_3664 : std_logic_vector(7 downto 0);
    signal wb27_3678 : std_logic_vector(7 downto 0);
    signal wb28_3692 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_3365_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3365_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3365_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3365_resized_base_address <= "00000000000000";
    array_obj_ref_3375_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3375_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3375_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3375_resized_base_address <= "00000000000000";
    konst_3277_wire_constant <= "0000000000000001";
    konst_3289_wire_constant <= "0000000000000001";
    konst_3291_wire_constant <= "0000000000000001";
    konst_3297_wire_constant <= "0000000000000001";
    konst_3300_wire_constant <= "0000000000000010";
    konst_3309_wire_constant <= "0000000000000001";
    konst_3362_wire_constant <= "00000000000000000000000000000011";
    konst_3372_wire_constant <= "00000000000000000000000000000011";
    konst_3471_wire_constant <= "000";
    konst_3485_wire_constant <= "001";
    konst_3499_wire_constant <= "010";
    konst_3513_wire_constant <= "011";
    konst_3527_wire_constant <= "100";
    konst_3541_wire_constant <= "101";
    konst_3555_wire_constant <= "110";
    konst_3569_wire_constant <= "111";
    konst_3583_wire_constant <= "000";
    konst_3597_wire_constant <= "001";
    konst_3611_wire_constant <= "010";
    konst_3625_wire_constant <= "011";
    konst_3639_wire_constant <= "100";
    konst_3653_wire_constant <= "101";
    konst_3667_wire_constant <= "110";
    konst_3681_wire_constant <= "111";
    konst_3737_wire_constant <= "0000000000000001";
    konst_3751_wire_constant <= "00000001";
    ptr_deref_3380_word_offset_0 <= "00000000000000";
    ptr_deref_3384_word_offset_0 <= "00000000000000";
    ptr_deref_3697_word_offset_0 <= "00000000000000";
    ptr_deref_3718_word_offset_0 <= "00000000000000";
    type_cast_3247_wire_constant <= "00000000000000000000000000000000";
    type_cast_3257_wire_constant <= "0000000000000000";
    type_cast_3262_wire_constant <= "0000000000000001";
    type_cast_3267_wire_constant <= "0000000000000001";
    phi_stmt_3244: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3247_wire_constant & n_address1_3343_3248_buffered;
      req <= phi_stmt_3244_req_0 & phi_stmt_3244_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3244",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3244_ack_0,
          idata => idata,
          odata => address1_3244,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3244
    phi_stmt_3249: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3252_wire & n_address2_3357_3253_buffered;
      req <= phi_stmt_3249_req_0 & phi_stmt_3249_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3249",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3249_ack_0,
          idata => idata,
          odata => address2_3249,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3249
    phi_stmt_3254: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3257_wire_constant & n_chl_3313_3258_buffered;
      req <= phi_stmt_3254_req_0 & phi_stmt_3254_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3254",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3254_ack_0,
          idata => idata,
          odata => chl_3254,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3254
    phi_stmt_3259: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3262_wire_constant & n_col_3294_3263_buffered;
      req <= phi_stmt_3259_req_0 & phi_stmt_3259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3259",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3259_ack_0,
          idata => idata,
          odata => col_3259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3259
    phi_stmt_3264: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3267_wire_constant & n_row_3305_3268_buffered;
      req <= phi_stmt_3264_req_0 & phi_stmt_3264_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3264",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3264_ack_0,
          idata => idata,
          odata => row_3264,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3264
    -- flow-through select operator MUX_3293_inst
    n_col_3294 <= konst_3289_wire_constant when (row_change_3274(0) /=  '0') else ADD_u16_u16_3292_wire;
    -- flow-through select operator MUX_3303_inst
    MUX_3303_wire <= ADD_u16_u16_3301_wire when (row_change_3274(0) /=  '0') else row_3264;
    -- flow-through select operator MUX_3304_inst
    n_row_3305 <= konst_3297_wire_constant when (chl_change_3286(0) /=  '0') else MUX_3303_wire;
    -- flow-through select operator MUX_3312_inst
    n_chl_3313 <= ADD_u16_u16_3310_wire when (chl_change_3286(0) /=  '0') else chl_3254;
    -- flow-through select operator MUX_3341_inst
    MUX_3341_wire <= ADD_u32_u32_3339_wire when (row_change_3274(0) /=  '0') else tmp1_3322;
    -- flow-through select operator MUX_3342_inst
    n_address1_3343 <= type_cast_3335_wire when (chl_change_3286(0) /=  '0') else MUX_3341_wire;
    -- flow-through select operator MUX_3355_inst
    MUX_3355_wire <= ADD_u32_u32_3353_wire when (row_change_3274(0) /=  '0') else tmp2_3331;
    -- flow-through select operator MUX_3356_inst
    n_address2_3357 <= ADD_u32_u32_3349_wire when (chl_change_3286(0) /=  '0') else MUX_3355_wire;
    -- flow-through select operator MUX_3481_inst
    wb11_3482 <= output_data1_3383_delayed_13_0_3476 when (EQ_u3_u1_3382_3382_delayed_14_0_3473(0) /=  '0') else w11_3400;
    -- flow-through select operator MUX_3495_inst
    wb12_3496 <= output_data1_3391_delayed_13_0_3490 when (EQ_u3_u1_3390_3390_delayed_14_0_3487(0) /=  '0') else w12_3404;
    -- flow-through select operator MUX_3509_inst
    wb13_3510 <= output_data1_3399_delayed_13_0_3504 when (EQ_u3_u1_3398_3398_delayed_14_0_3501(0) /=  '0') else w13_3408;
    -- flow-through select operator MUX_3523_inst
    wb14_3524 <= output_data1_3407_delayed_13_0_3518 when (EQ_u3_u1_3406_3406_delayed_14_0_3515(0) /=  '0') else w14_3412;
    -- flow-through select operator MUX_3537_inst
    wb15_3538 <= output_data1_3415_delayed_13_0_3532 when (EQ_u3_u1_3414_3414_delayed_14_0_3529(0) /=  '0') else w15_3416;
    -- flow-through select operator MUX_3551_inst
    wb16_3552 <= output_data1_3423_delayed_13_0_3546 when (EQ_u3_u1_3422_3422_delayed_14_0_3543(0) /=  '0') else w16_3420;
    -- flow-through select operator MUX_3565_inst
    wb17_3566 <= output_data1_3431_delayed_13_0_3560 when (EQ_u3_u1_3430_3430_delayed_14_0_3557(0) /=  '0') else w17_3424;
    -- flow-through select operator MUX_3579_inst
    wb18_3580 <= output_data1_3439_delayed_13_0_3574 when (EQ_u3_u1_3438_3438_delayed_14_0_3571(0) /=  '0') else w18_3428;
    -- flow-through select operator MUX_3593_inst
    wb21_3594 <= output_data2_3447_delayed_13_0_3588 when (EQ_u3_u1_3446_3446_delayed_14_0_3585(0) /=  '0') else w21_3432;
    -- flow-through select operator MUX_3607_inst
    wb22_3608 <= output_data2_3455_delayed_13_0_3602 when (EQ_u3_u1_3454_3454_delayed_14_0_3599(0) /=  '0') else w22_3436;
    -- flow-through select operator MUX_3621_inst
    wb23_3622 <= output_data2_3463_delayed_13_0_3616 when (EQ_u3_u1_3462_3462_delayed_14_0_3613(0) /=  '0') else w23_3440;
    -- flow-through select operator MUX_3635_inst
    wb24_3636 <= output_data2_3471_delayed_13_0_3630 when (EQ_u3_u1_3470_3470_delayed_14_0_3627(0) /=  '0') else w24_3444;
    -- flow-through select operator MUX_3649_inst
    wb25_3650 <= output_data2_3479_delayed_13_0_3644 when (EQ_u3_u1_3478_3478_delayed_14_0_3641(0) /=  '0') else w25_3448;
    -- flow-through select operator MUX_3663_inst
    wb26_3664 <= output_data2_3487_delayed_13_0_3658 when (EQ_u3_u1_3486_3486_delayed_14_0_3655(0) /=  '0') else w26_3452;
    -- flow-through select operator MUX_3677_inst
    wb27_3678 <= output_data2_3495_delayed_13_0_3672 when (EQ_u3_u1_3494_3494_delayed_14_0_3669(0) /=  '0') else w27_3456;
    -- flow-through select operator MUX_3691_inst
    wb28_3692 <= output_data2_3503_delayed_13_0_3686 when (EQ_u3_u1_3502_3502_delayed_14_0_3683(0) /=  '0') else w28_3460;
    slice_3391_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3391_inst_req_0;
      slice_3391_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3391_inst_req_1;
      slice_3391_inst_ack_1<= update_ack(0);
      slice_3391_inst: SliceSplitProtocol generic map(name => "slice_3391_inst", in_data_width => 16, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => output_data_read_3388, dout => output_data1_3392, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3395_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3395_inst_req_0;
      slice_3395_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3395_inst_req_1;
      slice_3395_inst_ack_1<= update_ack(0);
      slice_3395_inst: SliceSplitProtocol generic map(name => "slice_3395_inst", in_data_width => 16, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => output_data_read_3388, dout => output_data2_3396, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3399_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3399_inst_req_0;
      slice_3399_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3399_inst_req_1;
      slice_3399_inst_ack_1<= update_ack(0);
      slice_3399_inst: SliceSplitProtocol generic map(name => "slice_3399_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w11_3400, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3403_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3403_inst_req_0;
      slice_3403_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3403_inst_req_1;
      slice_3403_inst_ack_1<= update_ack(0);
      slice_3403_inst: SliceSplitProtocol generic map(name => "slice_3403_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w12_3404, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3407_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3407_inst_req_0;
      slice_3407_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3407_inst_req_1;
      slice_3407_inst_ack_1<= update_ack(0);
      slice_3407_inst: SliceSplitProtocol generic map(name => "slice_3407_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w13_3408, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3411_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3411_inst_req_0;
      slice_3411_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3411_inst_req_1;
      slice_3411_inst_ack_1<= update_ack(0);
      slice_3411_inst: SliceSplitProtocol generic map(name => "slice_3411_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w14_3412, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3415_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3415_inst_req_0;
      slice_3415_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3415_inst_req_1;
      slice_3415_inst_ack_1<= update_ack(0);
      slice_3415_inst: SliceSplitProtocol generic map(name => "slice_3415_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w15_3416, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3419_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3419_inst_req_0;
      slice_3419_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3419_inst_req_1;
      slice_3419_inst_ack_1<= update_ack(0);
      slice_3419_inst: SliceSplitProtocol generic map(name => "slice_3419_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w16_3420, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3423_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3423_inst_req_0;
      slice_3423_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3423_inst_req_1;
      slice_3423_inst_ack_1<= update_ack(0);
      slice_3423_inst: SliceSplitProtocol generic map(name => "slice_3423_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w17_3424, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3427_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3427_inst_req_0;
      slice_3427_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3427_inst_req_1;
      slice_3427_inst_ack_1<= update_ack(0);
      slice_3427_inst: SliceSplitProtocol generic map(name => "slice_3427_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val1_3381, dout => w18_3428, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3431_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3431_inst_req_0;
      slice_3431_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3431_inst_req_1;
      slice_3431_inst_ack_1<= update_ack(0);
      slice_3431_inst: SliceSplitProtocol generic map(name => "slice_3431_inst", in_data_width => 64, high_index => 63, low_index => 56, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w21_3432, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3435_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3435_inst_req_0;
      slice_3435_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3435_inst_req_1;
      slice_3435_inst_ack_1<= update_ack(0);
      slice_3435_inst: SliceSplitProtocol generic map(name => "slice_3435_inst", in_data_width => 64, high_index => 55, low_index => 48, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w22_3436, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3439_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3439_inst_req_0;
      slice_3439_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3439_inst_req_1;
      slice_3439_inst_ack_1<= update_ack(0);
      slice_3439_inst: SliceSplitProtocol generic map(name => "slice_3439_inst", in_data_width => 64, high_index => 47, low_index => 40, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w23_3440, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3443_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3443_inst_req_0;
      slice_3443_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3443_inst_req_1;
      slice_3443_inst_ack_1<= update_ack(0);
      slice_3443_inst: SliceSplitProtocol generic map(name => "slice_3443_inst", in_data_width => 64, high_index => 39, low_index => 32, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w24_3444, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3447_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3447_inst_req_0;
      slice_3447_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3447_inst_req_1;
      slice_3447_inst_ack_1<= update_ack(0);
      slice_3447_inst: SliceSplitProtocol generic map(name => "slice_3447_inst", in_data_width => 64, high_index => 31, low_index => 24, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w25_3448, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3451_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3451_inst_req_0;
      slice_3451_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3451_inst_req_1;
      slice_3451_inst_ack_1<= update_ack(0);
      slice_3451_inst: SliceSplitProtocol generic map(name => "slice_3451_inst", in_data_width => 64, high_index => 23, low_index => 16, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w26_3452, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3455_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3455_inst_req_0;
      slice_3455_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3455_inst_req_1;
      slice_3455_inst_ack_1<= update_ack(0);
      slice_3455_inst: SliceSplitProtocol generic map(name => "slice_3455_inst", in_data_width => 64, high_index => 15, low_index => 8, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w27_3456, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    slice_3459_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_3459_inst_req_0;
      slice_3459_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_3459_inst_req_1;
      slice_3459_inst_ack_1<= update_ack(0);
      slice_3459_inst: SliceSplitProtocol generic map(name => "slice_3459_inst", in_data_width => 64, high_index => 7, low_index => 0, buffering => 1, flow_through => false,  full_rate => true) -- 
        port map( din => fetch_val2_3385, dout => w28_3460, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    W_fetch_addr1_3507_delayed_8_0_3693_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr1_3507_delayed_8_0_3693_inst_req_0;
      W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr1_3507_delayed_8_0_3693_inst_req_1;
      W_fetch_addr1_3507_delayed_8_0_3693_inst_ack_1<= rack(0);
      W_fetch_addr1_3507_delayed_8_0_3693_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr1_3507_delayed_8_0_3693_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr1_3367,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3507_delayed_8_0_3695,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_fetch_addr2_3525_delayed_8_0_3714_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_fetch_addr2_3525_delayed_8_0_3714_inst_req_0;
      W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_0<= wack(0);
      rreq(0) <= W_fetch_addr2_3525_delayed_8_0_3714_inst_req_1;
      W_fetch_addr2_3525_delayed_8_0_3714_inst_ack_1<= rack(0);
      W_fetch_addr2_3525_delayed_8_0_3714_inst : InterlockBuffer generic map ( -- 
        name => "W_fetch_addr2_3525_delayed_8_0_3714_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => fetch_addr2_3377,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3525_delayed_8_0_3716,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3383_delayed_13_0_3474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3383_delayed_13_0_3474_inst_req_0;
      W_output_data1_3383_delayed_13_0_3474_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3383_delayed_13_0_3474_inst_req_1;
      W_output_data1_3383_delayed_13_0_3474_inst_ack_1<= rack(0);
      W_output_data1_3383_delayed_13_0_3474_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3383_delayed_13_0_3474_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3383_delayed_13_0_3476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3391_delayed_13_0_3488_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3391_delayed_13_0_3488_inst_req_0;
      W_output_data1_3391_delayed_13_0_3488_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3391_delayed_13_0_3488_inst_req_1;
      W_output_data1_3391_delayed_13_0_3488_inst_ack_1<= rack(0);
      W_output_data1_3391_delayed_13_0_3488_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3391_delayed_13_0_3488_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3391_delayed_13_0_3490,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3399_delayed_13_0_3502_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3399_delayed_13_0_3502_inst_req_0;
      W_output_data1_3399_delayed_13_0_3502_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3399_delayed_13_0_3502_inst_req_1;
      W_output_data1_3399_delayed_13_0_3502_inst_ack_1<= rack(0);
      W_output_data1_3399_delayed_13_0_3502_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3399_delayed_13_0_3502_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3399_delayed_13_0_3504,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3407_delayed_13_0_3516_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3407_delayed_13_0_3516_inst_req_0;
      W_output_data1_3407_delayed_13_0_3516_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3407_delayed_13_0_3516_inst_req_1;
      W_output_data1_3407_delayed_13_0_3516_inst_ack_1<= rack(0);
      W_output_data1_3407_delayed_13_0_3516_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3407_delayed_13_0_3516_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3407_delayed_13_0_3518,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3415_delayed_13_0_3530_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3415_delayed_13_0_3530_inst_req_0;
      W_output_data1_3415_delayed_13_0_3530_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3415_delayed_13_0_3530_inst_req_1;
      W_output_data1_3415_delayed_13_0_3530_inst_ack_1<= rack(0);
      W_output_data1_3415_delayed_13_0_3530_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3415_delayed_13_0_3530_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3415_delayed_13_0_3532,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3423_delayed_13_0_3544_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3423_delayed_13_0_3544_inst_req_0;
      W_output_data1_3423_delayed_13_0_3544_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3423_delayed_13_0_3544_inst_req_1;
      W_output_data1_3423_delayed_13_0_3544_inst_ack_1<= rack(0);
      W_output_data1_3423_delayed_13_0_3544_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3423_delayed_13_0_3544_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3423_delayed_13_0_3546,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3431_delayed_13_0_3558_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3431_delayed_13_0_3558_inst_req_0;
      W_output_data1_3431_delayed_13_0_3558_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3431_delayed_13_0_3558_inst_req_1;
      W_output_data1_3431_delayed_13_0_3558_inst_ack_1<= rack(0);
      W_output_data1_3431_delayed_13_0_3558_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3431_delayed_13_0_3558_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3431_delayed_13_0_3560,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data1_3439_delayed_13_0_3572_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data1_3439_delayed_13_0_3572_inst_req_0;
      W_output_data1_3439_delayed_13_0_3572_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data1_3439_delayed_13_0_3572_inst_req_1;
      W_output_data1_3439_delayed_13_0_3572_inst_ack_1<= rack(0);
      W_output_data1_3439_delayed_13_0_3572_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data1_3439_delayed_13_0_3572_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data1_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data1_3439_delayed_13_0_3574,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3447_delayed_13_0_3586_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3447_delayed_13_0_3586_inst_req_0;
      W_output_data2_3447_delayed_13_0_3586_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3447_delayed_13_0_3586_inst_req_1;
      W_output_data2_3447_delayed_13_0_3586_inst_ack_1<= rack(0);
      W_output_data2_3447_delayed_13_0_3586_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3447_delayed_13_0_3586_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3447_delayed_13_0_3588,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3455_delayed_13_0_3600_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3455_delayed_13_0_3600_inst_req_0;
      W_output_data2_3455_delayed_13_0_3600_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3455_delayed_13_0_3600_inst_req_1;
      W_output_data2_3455_delayed_13_0_3600_inst_ack_1<= rack(0);
      W_output_data2_3455_delayed_13_0_3600_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3455_delayed_13_0_3600_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3455_delayed_13_0_3602,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3463_delayed_13_0_3614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3463_delayed_13_0_3614_inst_req_0;
      W_output_data2_3463_delayed_13_0_3614_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3463_delayed_13_0_3614_inst_req_1;
      W_output_data2_3463_delayed_13_0_3614_inst_ack_1<= rack(0);
      W_output_data2_3463_delayed_13_0_3614_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3463_delayed_13_0_3614_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3463_delayed_13_0_3616,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3471_delayed_13_0_3628_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3471_delayed_13_0_3628_inst_req_0;
      W_output_data2_3471_delayed_13_0_3628_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3471_delayed_13_0_3628_inst_req_1;
      W_output_data2_3471_delayed_13_0_3628_inst_ack_1<= rack(0);
      W_output_data2_3471_delayed_13_0_3628_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3471_delayed_13_0_3628_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3471_delayed_13_0_3630,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3479_delayed_13_0_3642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3479_delayed_13_0_3642_inst_req_0;
      W_output_data2_3479_delayed_13_0_3642_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3479_delayed_13_0_3642_inst_req_1;
      W_output_data2_3479_delayed_13_0_3642_inst_ack_1<= rack(0);
      W_output_data2_3479_delayed_13_0_3642_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3479_delayed_13_0_3642_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3479_delayed_13_0_3644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3487_delayed_13_0_3656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3487_delayed_13_0_3656_inst_req_0;
      W_output_data2_3487_delayed_13_0_3656_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3487_delayed_13_0_3656_inst_req_1;
      W_output_data2_3487_delayed_13_0_3656_inst_ack_1<= rack(0);
      W_output_data2_3487_delayed_13_0_3656_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3487_delayed_13_0_3656_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3487_delayed_13_0_3658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3495_delayed_13_0_3670_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3495_delayed_13_0_3670_inst_req_0;
      W_output_data2_3495_delayed_13_0_3670_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3495_delayed_13_0_3670_inst_req_1;
      W_output_data2_3495_delayed_13_0_3670_inst_ack_1<= rack(0);
      W_output_data2_3495_delayed_13_0_3670_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3495_delayed_13_0_3670_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3495_delayed_13_0_3672,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_output_data2_3503_delayed_13_0_3684_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_output_data2_3503_delayed_13_0_3684_inst_req_0;
      W_output_data2_3503_delayed_13_0_3684_inst_ack_0<= wack(0);
      rreq(0) <= W_output_data2_3503_delayed_13_0_3684_inst_req_1;
      W_output_data2_3503_delayed_13_0_3684_inst_ack_1<= rack(0);
      W_output_data2_3503_delayed_13_0_3684_inst : InterlockBuffer generic map ( -- 
        name => "W_output_data2_3503_delayed_13_0_3684_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => output_data2_3396,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => output_data2_3503_delayed_13_0_3686,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3366_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3366_final_reg_req_0;
      addr_of_3366_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3366_final_reg_req_1;
      addr_of_3366_final_reg_ack_1<= rack(0);
      addr_of_3366_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3366_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3365_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr1_3367,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3376_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3376_final_reg_req_0;
      addr_of_3376_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3376_final_reg_req_1;
      addr_of_3376_final_reg_ack_1<= rack(0);
      addr_of_3376_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3376_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3375_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => fetch_addr2_3377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address1_3343_3248_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address1_3343_3248_buf_req_0;
      n_address1_3343_3248_buf_ack_0<= wack(0);
      rreq(0) <= n_address1_3343_3248_buf_req_1;
      n_address1_3343_3248_buf_ack_1<= rack(0);
      n_address1_3343_3248_buf : InterlockBuffer generic map ( -- 
        name => "n_address1_3343_3248_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address1_3343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address1_3343_3248_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_address2_3357_3253_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_address2_3357_3253_buf_req_0;
      n_address2_3357_3253_buf_ack_0<= wack(0);
      rreq(0) <= n_address2_3357_3253_buf_req_1;
      n_address2_3357_3253_buf_ack_1<= rack(0);
      n_address2_3357_3253_buf : InterlockBuffer generic map ( -- 
        name => "n_address2_3357_3253_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_address2_3357,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_address2_3357_3253_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_chl_3313_3258_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_chl_3313_3258_buf_req_0;
      n_chl_3313_3258_buf_ack_0<= wack(0);
      rreq(0) <= n_chl_3313_3258_buf_req_1;
      n_chl_3313_3258_buf_ack_1<= rack(0);
      n_chl_3313_3258_buf : InterlockBuffer generic map ( -- 
        name => "n_chl_3313_3258_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_chl_3313,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_chl_3313_3258_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_col_3294_3263_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_col_3294_3263_buf_req_0;
      n_col_3294_3263_buf_ack_0<= wack(0);
      rreq(0) <= n_col_3294_3263_buf_req_1;
      n_col_3294_3263_buf_ack_1<= rack(0);
      n_col_3294_3263_buf : InterlockBuffer generic map ( -- 
        name => "n_col_3294_3263_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_col_3294,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_col_3294_3263_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_row_3305_3268_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_row_3305_3268_buf_req_0;
      n_row_3305_3268_buf_ack_0<= wack(0);
      rreq(0) <= n_row_3305_3268_buf_req_1;
      n_row_3305_3268_buf_ack_1<= rack(0);
      n_row_3305_3268_buf : InterlockBuffer generic map ( -- 
        name => "n_row_3305_3268_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_row_3305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_row_3305_3268_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3240_inst
    process(MUL_u16_u16_3239_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := MUL_u16_u16_3239_wire(15 downto 0);
      row_size_3241 <= tmp_var; -- 
    end process;
    type_cast_3252_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3252_inst_req_0;
      type_cast_3252_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3252_inst_req_1;
      type_cast_3252_inst_ack_1<= rack(0);
      type_cast_3252_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3252_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => row_size_3241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3252_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3316_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3316_inst_req_0;
      type_cast_3316_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3316_inst_req_1;
      type_cast_3316_inst_ack_1<= rack(0);
      type_cast_3316_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3316_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3233_3233_delayed_1_0_3317,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3325_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3325_inst_req_0;
      type_cast_3325_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3325_inst_req_1;
      type_cast_3325_inst_ack_1<= rack(0);
      type_cast_3325_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3325_inst",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => chl_out_3235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3239_3239_delayed_1_0_3326,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3335_inst
    process(n_chl_3313) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3313(15 downto 0);
      type_cast_3335_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3347_inst
    process(n_chl_3313) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := n_chl_3313(15 downto 0);
      type_cast_3347_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3364_inst
    process(LSHR_u32_u32_3363_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3363_wire(31 downto 0);
      type_cast_3364_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3374_inst
    process(LSHR_u32_u32_3373_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := LSHR_u32_u32_3373_wire(31 downto 0);
      type_cast_3374_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3463_inst
    process(address1_3244) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := address1_3244(2 downto 0);
      location1_3464 <= tmp_var; -- 
    end process;
    -- interlock type_cast_3467_inst
    process(address2_3249) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := address2_3249(2 downto 0);
      location2_3468 <= tmp_var; -- 
    end process;
    -- equivalence array_obj_ref_3365_index_1_rename
    process(type_cast_3364_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3364_resized;
      ov(13 downto 0) := iv;
      type_cast_3364_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3365_index_1_resize
    process(type_cast_3364_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3364_wire;
      ov := iv(13 downto 0);
      type_cast_3364_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3365_root_address_inst
    process(array_obj_ref_3365_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3365_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3365_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3375_index_1_rename
    process(type_cast_3374_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3374_resized;
      ov(13 downto 0) := iv;
      type_cast_3374_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3375_index_1_resize
    process(type_cast_3374_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_3374_wire;
      ov := iv(13 downto 0);
      type_cast_3374_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3375_root_address_inst
    process(array_obj_ref_3375_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3375_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3375_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3380_addr_0
    process(ptr_deref_3380_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3380_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3380_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3380_base_resize
    process(fetch_addr1_3367) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3367;
      ov := iv(13 downto 0);
      ptr_deref_3380_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3380_gather_scatter
    process(ptr_deref_3380_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3380_data_0;
      ov(63 downto 0) := iv;
      fetch_val1_3381 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3380_root_address_inst
    process(ptr_deref_3380_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3380_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3380_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3384_addr_0
    process(ptr_deref_3384_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3384_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3384_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3384_base_resize
    process(fetch_addr2_3377) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3377;
      ov := iv(13 downto 0);
      ptr_deref_3384_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3384_gather_scatter
    process(ptr_deref_3384_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3384_data_0;
      ov(63 downto 0) := iv;
      fetch_val2_3385 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3384_root_address_inst
    process(ptr_deref_3384_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3384_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3384_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3697_addr_0
    process(ptr_deref_3697_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3697_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3697_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3697_base_resize
    process(fetch_addr1_3507_delayed_8_0_3695) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr1_3507_delayed_8_0_3695;
      ov := iv(13 downto 0);
      ptr_deref_3697_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3697_gather_scatter
    process(CONCAT_u32_u64_3712_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3712_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3697_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3697_root_address_inst
    process(ptr_deref_3697_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3697_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3697_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3718_addr_0
    process(ptr_deref_3718_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3718_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3718_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3718_base_resize
    process(fetch_addr2_3525_delayed_8_0_3716) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := fetch_addr2_3525_delayed_8_0_3716;
      ov := iv(13 downto 0);
      ptr_deref_3718_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3718_gather_scatter
    process(CONCAT_u32_u64_3733_wire) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := CONCAT_u32_u64_3733_wire;
      ov(63 downto 0) := iv;
      ptr_deref_3718_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3718_root_address_inst
    process(ptr_deref_3718_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3718_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3718_root_address <= ov(13 downto 0);
      --
    end process;
    do_while_stmt_3242_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3747;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3242_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3242_branch_req_0,
          ack0 => do_while_stmt_3242_branch_ack_0,
          ack1 => do_while_stmt_3242_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3292_inst
    process(col_3259) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(col_3259, konst_3291_wire_constant, tmp_var);
      ADD_u16_u16_3292_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3301_inst
    process(row_3264) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(row_3264, konst_3300_wire_constant, tmp_var);
      ADD_u16_u16_3301_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3310_inst
    process(chl_3254) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(chl_3254, konst_3309_wire_constant, tmp_var);
      ADD_u16_u16_3310_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3321_inst
    process(address1_3244, type_cast_3233_3233_delayed_1_0_3317) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address1_3244, type_cast_3233_3233_delayed_1_0_3317, tmp_var);
      tmp1_3322 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3330_inst
    process(address2_3249, type_cast_3239_3239_delayed_1_0_3326) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(address2_3249, type_cast_3239_3239_delayed_1_0_3326, tmp_var);
      tmp2_3331 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3339_inst
    process(tmp1_3322, row_size_3241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp1_3322, row_size_3241, tmp_var);
      ADD_u32_u32_3339_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3349_inst
    process(type_cast_3347_wire, row_size_3241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(type_cast_3347_wire, row_size_3241, tmp_var);
      ADD_u32_u32_3349_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3353_inst
    process(tmp2_3331, row_size_3241) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp2_3331, row_size_3241, tmp_var);
      ADD_u32_u32_3353_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3285_inst
    process(row_change_3274, UGE_u16_u1_3284_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(row_change_3274, UGE_u16_u1_3284_wire, tmp_var);
      chl_change_3286 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3704_inst
    process(CONCAT_u8_u16_3700_wire, CONCAT_u8_u16_3703_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3700_wire, CONCAT_u8_u16_3703_wire, tmp_var);
      CONCAT_u16_u32_3704_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3711_inst
    process(CONCAT_u8_u16_3707_wire, CONCAT_u8_u16_3710_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3707_wire, CONCAT_u8_u16_3710_wire, tmp_var);
      CONCAT_u16_u32_3711_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3725_inst
    process(CONCAT_u8_u16_3721_wire, CONCAT_u8_u16_3724_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3721_wire, CONCAT_u8_u16_3724_wire, tmp_var);
      CONCAT_u16_u32_3725_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_3732_inst
    process(CONCAT_u8_u16_3728_wire, CONCAT_u8_u16_3731_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_3728_wire, CONCAT_u8_u16_3731_wire, tmp_var);
      CONCAT_u16_u32_3732_wire <= tmp_var; --
    end process;
    -- shared split operator group (13) : CONCAT_u32_u64_3712_inst 
    ApConcat_group_13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3704_wire & CONCAT_u16_u32_3711_wire;
      CONCAT_u32_u64_3712_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3712_inst_req_0;
      CONCAT_u32_u64_3712_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3712_inst_req_1;
      CONCAT_u32_u64_3712_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_13_gI: SplitGuardInterface generic map(name => "ApConcat_group_13_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_13",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : CONCAT_u32_u64_3733_inst 
    ApConcat_group_14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u32_3725_wire & CONCAT_u16_u32_3732_wire;
      CONCAT_u32_u64_3733_wire <= data_out(63 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u32_u64_3733_inst_req_0;
      CONCAT_u32_u64_3733_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u32_u64_3733_inst_req_1;
      CONCAT_u32_u64_3733_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_14_gI: SplitGuardInterface generic map(name => "ApConcat_group_14_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_14",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- binary operator CONCAT_u8_u16_3700_inst
    process(wb11_3482, wb12_3496) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb11_3482, wb12_3496, tmp_var);
      CONCAT_u8_u16_3700_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3703_inst
    process(wb13_3510, wb14_3524) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb13_3510, wb14_3524, tmp_var);
      CONCAT_u8_u16_3703_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3707_inst
    process(wb15_3538, wb16_3552) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb15_3538, wb16_3552, tmp_var);
      CONCAT_u8_u16_3707_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3710_inst
    process(wb17_3566, wb18_3580) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb17_3566, wb18_3580, tmp_var);
      CONCAT_u8_u16_3710_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3721_inst
    process(wb21_3594, wb22_3608) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb21_3594, wb22_3608, tmp_var);
      CONCAT_u8_u16_3721_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3724_inst
    process(wb23_3622, wb24_3636) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb23_3622, wb24_3636, tmp_var);
      CONCAT_u8_u16_3724_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3728_inst
    process(wb25_3650, wb26_3664) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb25_3650, wb26_3664, tmp_var);
      CONCAT_u8_u16_3728_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_3731_inst
    process(wb27_3678, wb28_3692) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(wb27_3678, wb28_3692, tmp_var);
      CONCAT_u8_u16_3731_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u16_u1_3273_inst
    process(col_3259, cb_3232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(col_3259, cb_3232, tmp_var);
      row_change_3274 <= tmp_var; --
    end process;
    -- shared split operator group (24) : EQ_u3_u1_3472_inst 
    ApIntEq_group_24: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3382_3382_delayed_14_0_3473 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3472_inst_req_0;
      EQ_u3_u1_3472_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3472_inst_req_1;
      EQ_u3_u1_3472_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_24_gI: SplitGuardInterface generic map(name => "ApIntEq_group_24_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_24",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : EQ_u3_u1_3486_inst 
    ApIntEq_group_25: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3390_3390_delayed_14_0_3487 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3486_inst_req_0;
      EQ_u3_u1_3486_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3486_inst_req_1;
      EQ_u3_u1_3486_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_25_gI: SplitGuardInterface generic map(name => "ApIntEq_group_25_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_25",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "001",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : EQ_u3_u1_3500_inst 
    ApIntEq_group_26: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3398_3398_delayed_14_0_3501 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3500_inst_req_0;
      EQ_u3_u1_3500_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3500_inst_req_1;
      EQ_u3_u1_3500_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_26_gI: SplitGuardInterface generic map(name => "ApIntEq_group_26_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_26",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "010",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : EQ_u3_u1_3514_inst 
    ApIntEq_group_27: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3406_3406_delayed_14_0_3515 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3514_inst_req_0;
      EQ_u3_u1_3514_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3514_inst_req_1;
      EQ_u3_u1_3514_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_27_gI: SplitGuardInterface generic map(name => "ApIntEq_group_27_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_27",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "011",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : EQ_u3_u1_3528_inst 
    ApIntEq_group_28: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3414_3414_delayed_14_0_3529 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3528_inst_req_0;
      EQ_u3_u1_3528_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3528_inst_req_1;
      EQ_u3_u1_3528_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_28_gI: SplitGuardInterface generic map(name => "ApIntEq_group_28_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_28",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : EQ_u3_u1_3542_inst 
    ApIntEq_group_29: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3422_3422_delayed_14_0_3543 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3542_inst_req_0;
      EQ_u3_u1_3542_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3542_inst_req_1;
      EQ_u3_u1_3542_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_29_gI: SplitGuardInterface generic map(name => "ApIntEq_group_29_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_29",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "101",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : EQ_u3_u1_3556_inst 
    ApIntEq_group_30: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3430_3430_delayed_14_0_3557 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3556_inst_req_0;
      EQ_u3_u1_3556_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3556_inst_req_1;
      EQ_u3_u1_3556_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_30_gI: SplitGuardInterface generic map(name => "ApIntEq_group_30_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_30",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "110",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : EQ_u3_u1_3570_inst 
    ApIntEq_group_31: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location1_3464;
      EQ_u3_u1_3438_3438_delayed_14_0_3571 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3570_inst_req_0;
      EQ_u3_u1_3570_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3570_inst_req_1;
      EQ_u3_u1_3570_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_31_gI: SplitGuardInterface generic map(name => "ApIntEq_group_31_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_31",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "111",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : EQ_u3_u1_3584_inst 
    ApIntEq_group_32: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3446_3446_delayed_14_0_3585 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3584_inst_req_0;
      EQ_u3_u1_3584_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3584_inst_req_1;
      EQ_u3_u1_3584_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_32_gI: SplitGuardInterface generic map(name => "ApIntEq_group_32_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_32",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "000",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : EQ_u3_u1_3598_inst 
    ApIntEq_group_33: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3454_3454_delayed_14_0_3599 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3598_inst_req_0;
      EQ_u3_u1_3598_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3598_inst_req_1;
      EQ_u3_u1_3598_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_33_gI: SplitGuardInterface generic map(name => "ApIntEq_group_33_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_33",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "001",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : EQ_u3_u1_3612_inst 
    ApIntEq_group_34: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3462_3462_delayed_14_0_3613 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3612_inst_req_0;
      EQ_u3_u1_3612_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3612_inst_req_1;
      EQ_u3_u1_3612_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_34_gI: SplitGuardInterface generic map(name => "ApIntEq_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "010",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : EQ_u3_u1_3626_inst 
    ApIntEq_group_35: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3470_3470_delayed_14_0_3627 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3626_inst_req_0;
      EQ_u3_u1_3626_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3626_inst_req_1;
      EQ_u3_u1_3626_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_35_gI: SplitGuardInterface generic map(name => "ApIntEq_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "011",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : EQ_u3_u1_3640_inst 
    ApIntEq_group_36: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3478_3478_delayed_14_0_3641 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3640_inst_req_0;
      EQ_u3_u1_3640_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3640_inst_req_1;
      EQ_u3_u1_3640_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_36_gI: SplitGuardInterface generic map(name => "ApIntEq_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "100",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : EQ_u3_u1_3654_inst 
    ApIntEq_group_37: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3486_3486_delayed_14_0_3655 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3654_inst_req_0;
      EQ_u3_u1_3654_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3654_inst_req_1;
      EQ_u3_u1_3654_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_37_gI: SplitGuardInterface generic map(name => "ApIntEq_group_37_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_37",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "101",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : EQ_u3_u1_3668_inst 
    ApIntEq_group_38: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3494_3494_delayed_14_0_3669 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3668_inst_req_0;
      EQ_u3_u1_3668_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3668_inst_req_1;
      EQ_u3_u1_3668_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_38_gI: SplitGuardInterface generic map(name => "ApIntEq_group_38_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_38",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "110",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : EQ_u3_u1_3682_inst 
    ApIntEq_group_39: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= location2_3468;
      EQ_u3_u1_3502_3502_delayed_14_0_3683 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u3_u1_3682_inst_req_0;
      EQ_u3_u1_3682_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u3_u1_3682_inst_req_1;
      EQ_u3_u1_3682_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_39_gI: SplitGuardInterface generic map(name => "ApIntEq_group_39_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_39",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 3,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "111",
          constant_width => 3,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- binary operator LSHR_u32_u32_3363_inst
    process(address1_3244) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address1_3244, konst_3362_wire_constant, tmp_var);
      LSHR_u32_u32_3363_wire <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3373_inst
    process(address2_3249) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(address2_3249, konst_3372_wire_constant, tmp_var);
      LSHR_u32_u32_3373_wire <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3239_inst
    process(chl_out_3235, cb_3232) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(chl_out_3235, cb_3232, tmp_var);
      MUL_u16_u16_3239_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3745_inst
    process(chl_change_3286) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", chl_change_3286, tmp_var);
      NOT_u1_u1_3745_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3746_inst
    process(ULT_u16_u1_3743_wire, NOT_u1_u1_3745_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(ULT_u16_u1_3743_wire, NOT_u1_u1_3745_wire, tmp_var);
      continue_flag_3747 <= tmp_var; --
    end process;
    -- shared split operator group (45) : SUB_u16_u16_3278_inst 
    ApIntSub_group_45: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= rb_3229;
      SUB_u16_u16_3199_3199_delayed_1_0_3279 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3278_inst_req_0;
      SUB_u16_u16_3278_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3278_inst_req_1;
      SUB_u16_u16_3278_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_45_gI: SplitGuardInterface generic map(name => "ApIntSub_group_45_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_45",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : SUB_u16_u16_3738_inst 
    ApIntSub_group_46: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= chl_out_3235;
      SUB_u16_u16_3547_3547_delayed_1_0_3739 <= data_out(15 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u16_u16_3738_inst_req_0;
      SUB_u16_u16_3738_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u16_u16_3738_inst_req_1;
      SUB_u16_u16_3738_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_46_gI: SplitGuardInterface generic map(name => "ApIntSub_group_46_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_46",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- binary operator UGE_u16_u1_3284_inst
    process(row_3264, SUB_u16_u16_3199_3199_delayed_1_0_3279) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(row_3264, SUB_u16_u16_3199_3199_delayed_1_0_3279, tmp_var);
      UGE_u16_u1_3284_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u16_u1_3743_inst
    process(chl_3254, SUB_u16_u16_3547_3547_delayed_1_0_3739) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(chl_3254, SUB_u16_u16_3547_3547_delayed_1_0_3739, tmp_var);
      ULT_u16_u1_3743_wire <= tmp_var; --
    end process;
    -- shared split operator group (49) : array_obj_ref_3365_index_offset 
    ApIntAdd_group_49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3364_scaled;
      array_obj_ref_3365_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3365_index_offset_req_0;
      array_obj_ref_3365_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3365_index_offset_req_1;
      array_obj_ref_3365_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_49_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_49_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_49",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : array_obj_ref_3375_index_offset 
    ApIntAdd_group_50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= type_cast_3374_scaled;
      array_obj_ref_3375_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3375_index_offset_req_0;
      array_obj_ref_3375_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3375_index_offset_req_1;
      array_obj_ref_3375_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_50_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_50_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_50",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 2,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared load operator group (0) : ptr_deref_3384_load_0 ptr_deref_3380_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3384_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3380_load_0_req_0;
      ptr_deref_3384_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3380_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3384_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3380_load_0_req_1;
      ptr_deref_3384_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3380_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3384_word_address_0 & ptr_deref_3380_word_address_0;
      ptr_deref_3384_data_0 <= data_out(127 downto 64);
      ptr_deref_3380_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 14,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(13 downto 0),
          mtag => memory_space_0_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(63 downto 0),
          mtag => memory_space_0_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_3697_store_0 ptr_deref_3718_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(27 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 15, 0 => 15);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 6, 1 => 6);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_3697_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_3718_store_0_req_0;
      ptr_deref_3697_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_3718_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_3697_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_3718_store_0_req_1;
      ptr_deref_3697_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_3718_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup0_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_0", num_slots => 2) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup0_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup0_accessRegulator_1", num_slots => 2) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3697_word_address_0 & ptr_deref_3718_word_address_0;
      data_in <= ptr_deref_3697_data_0 & ptr_deref_3718_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 17,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(13 downto 0),
          mdata => memory_space_0_sr_data(63 downto 0),
          mtag => memory_space_0_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_output_pipe_3234_inst RPIPE_output_pipe_3231_inst RPIPE_output_pipe_3228_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(47 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 2 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= RPIPE_output_pipe_3234_inst_req_0;
      reqL_unguarded(1) <= RPIPE_output_pipe_3231_inst_req_0;
      reqL_unguarded(0) <= RPIPE_output_pipe_3228_inst_req_0;
      RPIPE_output_pipe_3234_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_output_pipe_3231_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_output_pipe_3228_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= RPIPE_output_pipe_3234_inst_req_1;
      reqR_unguarded(1) <= RPIPE_output_pipe_3231_inst_req_1;
      reqR_unguarded(0) <= RPIPE_output_pipe_3228_inst_req_1;
      RPIPE_output_pipe_3234_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_output_pipe_3231_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_output_pipe_3228_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      chl_out_3235 <= data_out(47 downto 32);
      cb_3232 <= data_out(31 downto 16);
      rb_3229 <= data_out(15 downto 0);
      output_pipe_read_0_gI: SplitGuardInterface generic map(name => "output_pipe_read_0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_0: InputPortRevised -- 
        generic map ( name => "output_pipe_read_0", data_width => 16,  num_reqs => 3,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(1),
          oack => output_pipe_pipe_read_ack(1),
          odata => output_pipe_pipe_read_data(31 downto 16),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_output_pipe_3387_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_output_pipe_3387_inst_req_0;
      RPIPE_output_pipe_3387_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_output_pipe_3387_inst_req_1;
      RPIPE_output_pipe_3387_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      output_data_read_3388 <= data_out(15 downto 0);
      output_pipe_read_1_gI: SplitGuardInterface generic map(name => "output_pipe_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      output_pipe_read_1: InputPortRevised -- 
        generic map ( name => "output_pipe_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => output_pipe_pipe_read_req(0),
          oack => output_pipe_pipe_read_ack(0),
          odata => output_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : WPIPE_input_done_pipe_3750_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_input_done_pipe_3750_inst_req_0;
      WPIPE_input_done_pipe_3750_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_input_done_pipe_3750_inst_req_1;
      WPIPE_input_done_pipe_3750_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_3751_wire_constant;
      input_done_pipe_write_0_gI: SplitGuardInterface generic map(name => "input_done_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      input_done_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "input_done_pipe", data_width => 8, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => input_done_pipe_pipe_write_req(0),
          oack => input_done_pipe_pipe_write_ack(0),
          odata => input_done_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendModule_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timer is -- 
  generic (tag_length : integer); 
  port ( -- 
    T : out  std_logic_vector(63 downto 0);
    timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
    timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timer;
architecture timer_arch of timer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal T_buffer :  std_logic_vector(63 downto 0);
  signal T_update_enable: Boolean;
  signal timer_CP_1315_start: Boolean;
  signal timer_CP_1315_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_timer_resp_408_inst_req_0 : boolean;
  signal WPIPE_timer_req_403_inst_ack_1 : boolean;
  signal WPIPE_timer_req_403_inst_req_1 : boolean;
  signal WPIPE_timer_req_403_inst_req_0 : boolean;
  signal WPIPE_timer_req_403_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_408_inst_ack_0 : boolean;
  signal RPIPE_timer_resp_408_inst_req_1 : boolean;
  signal RPIPE_timer_resp_408_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timer_CP_1315_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= T_buffer;
  T <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1315_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timer_CP_1315_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timer_CP_1315_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timer_CP_1315: Block -- control-path 
    signal timer_CP_1315_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    timer_CP_1315_elements(0) <= timer_CP_1315_start;
    timer_CP_1315_symbol <= timer_CP_1315_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_sample_start_
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Sample/rr
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_sample_start_
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/$entry
      -- CP-element group 0: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Sample/req
      -- CP-element group 0: 	 $entry
      -- 
    rr_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1315_elements(0), ack => RPIPE_timer_resp_408_inst_req_0); -- 
    req_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1315_elements(0), ack => WPIPE_timer_req_403_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_sample_completed_
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Update/req
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Update/$entry
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_update_start_
      -- CP-element group 1: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Sample/ack
      -- 
    ack_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_403_inst_ack_0, ack => timer_CP_1315_elements(1)); -- 
    req_1333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1315_elements(1), ack => WPIPE_timer_req_403_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_update_completed_
      -- CP-element group 2: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Update/ack
      -- CP-element group 2: 	 assign_stmt_406_to_assign_stmt_409/WPIPE_timer_req_403_Update/$exit
      -- 
    ack_1334_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_req_403_inst_ack_1, ack => timer_CP_1315_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_update_start_
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_sample_completed_
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Sample/ra
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Update/$entry
      -- CP-element group 3: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Update/cr
      -- 
    ra_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_408_inst_ack_0, ack => timer_CP_1315_elements(3)); -- 
    cr_1347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timer_CP_1315_elements(3), ack => RPIPE_timer_resp_408_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_update_completed_
      -- CP-element group 4: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Update/$exit
      -- CP-element group 4: 	 assign_stmt_406_to_assign_stmt_409/RPIPE_timer_resp_408_Update/ca
      -- 
    ca_1348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_resp_408_inst_ack_1, ack => timer_CP_1315_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_406_to_assign_stmt_409/$exit
      -- 
    timer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 24) := "timer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timer_CP_1315_elements(4) & timer_CP_1315_elements(2);
      gj_timer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timer_CP_1315_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal type_cast_405_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_405_wire_constant <= "1";
    -- shared inport operator group (0) : RPIPE_timer_resp_408_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_resp_408_inst_req_0;
      RPIPE_timer_resp_408_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_resp_408_inst_req_1;
      RPIPE_timer_resp_408_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      T_buffer <= data_out(63 downto 0);
      timer_resp_read_0_gI: SplitGuardInterface generic map(name => "timer_resp_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_resp_read_0: InputPortRevised -- 
        generic map ( name => "timer_resp_read_0", data_width => 64,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_resp_pipe_read_req(0),
          oack => timer_resp_pipe_read_ack(0),
          odata => timer_resp_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_req_403_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_req_403_inst_req_0;
      WPIPE_timer_req_403_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_req_403_inst_req_1;
      WPIPE_timer_req_403_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_405_wire_constant;
      timer_req_write_0_gI: SplitGuardInterface generic map(name => "timer_req_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_req_write_0: OutputPortRevised -- 
        generic map ( name => "timer_req", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_req_pipe_write_req(0),
          oack => timer_req_pipe_write_ack(0),
          odata => timer_req_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity timerDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
    timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
    timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
    timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
    timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity timerDaemon;
architecture timerDaemon_arch of timerDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal timerDaemon_CP_9188_start: Boolean;
  signal timerDaemon_CP_9188_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_timer_resp_4061_inst_req_0 : boolean;
  signal WPIPE_timer_resp_4061_inst_ack_0 : boolean;
  signal do_while_stmt_4044_branch_ack_0 : boolean;
  signal do_while_stmt_4044_branch_ack_1 : boolean;
  signal WPIPE_timer_resp_4061_inst_req_1 : boolean;
  signal WPIPE_timer_resp_4061_inst_ack_1 : boolean;
  signal do_while_stmt_4044_branch_req_0 : boolean;
  signal phi_stmt_4046_req_0 : boolean;
  signal phi_stmt_4046_req_1 : boolean;
  signal phi_stmt_4046_ack_0 : boolean;
  signal nCOUNTER_4059_4048_buf_req_0 : boolean;
  signal nCOUNTER_4059_4048_buf_ack_0 : boolean;
  signal nCOUNTER_4059_4048_buf_req_1 : boolean;
  signal nCOUNTER_4059_4048_buf_ack_1 : boolean;
  signal RPIPE_timer_req_4053_inst_req_0 : boolean;
  signal RPIPE_timer_req_4053_inst_ack_0 : boolean;
  signal RPIPE_timer_req_4053_inst_req_1 : boolean;
  signal RPIPE_timer_req_4053_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "timerDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  timerDaemon_CP_9188_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "timerDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_9188_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= timerDaemon_CP_9188_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= timerDaemon_CP_9188_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  timerDaemon_CP_9188: Block -- control-path 
    signal timerDaemon_CP_9188_elements: BooleanArray(44 downto 0);
    -- 
  begin -- 
    timerDaemon_CP_9188_elements(0) <= timerDaemon_CP_9188_start;
    timerDaemon_CP_9188_symbol <= timerDaemon_CP_9188_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_4043/$entry
      -- CP-element group 0: 	 branch_block_stmt_4043/branch_block_stmt_4043__entry__
      -- CP-element group 0: 	 branch_block_stmt_4043/do_while_stmt_4044__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	44 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_4043/$exit
      -- CP-element group 1: 	 branch_block_stmt_4043/branch_block_stmt_4043__exit__
      -- CP-element group 1: 	 branch_block_stmt_4043/do_while_stmt_4044__exit__
      -- 
    timerDaemon_CP_9188_elements(1) <= timerDaemon_CP_9188_elements(44);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_4043/do_while_stmt_4044/$entry
      -- CP-element group 2: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044__entry__
      -- 
    timerDaemon_CP_9188_elements(2) <= timerDaemon_CP_9188_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	44 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044__exit__
      -- 
    -- Element group timerDaemon_CP_9188_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_back
      -- 
    -- Element group timerDaemon_CP_9188_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	42 
    -- CP-element group 5: 	43 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_4043/do_while_stmt_4044/condition_done
      -- 
    timerDaemon_CP_9188_elements(5) <= timerDaemon_CP_9188_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	41 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_body_done
      -- 
    timerDaemon_CP_9188_elements(6) <= timerDaemon_CP_9188_elements(41);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/back_edge_to_loop_body
      -- 
    timerDaemon_CP_9188_elements(7) <= timerDaemon_CP_9188_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/first_time_through_loop_body
      -- 
    timerDaemon_CP_9188_elements(8) <= timerDaemon_CP_9188_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	32 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4051_sample_start_
      -- 
    -- Element group timerDaemon_CP_9188_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	40 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/condition_evaluated
      -- 
    condition_evaluated_9212_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_9212_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(10), ack => do_while_stmt_4044_branch_req_0); -- 
    timerDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(40) & timerDaemon_CP_9188_elements(14);
      gj_timerDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	33 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_sample_start__ps
      -- 
    timerDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(15) & timerDaemon_CP_9188_elements(9) & timerDaemon_CP_9188_elements(14);
      gj_timerDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	35 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	41 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4051_sample_completed_
      -- 
    timerDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(35) & timerDaemon_CP_9188_elements(17);
      gj_timerDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	32 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	34 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_update_start__ps
      -- 
    timerDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(32) & timerDaemon_CP_9188_elements(16);
      gj_timerDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	36 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/aggregated_phi_update_ack
      -- 
    timerDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(36) & timerDaemon_CP_9188_elements(18);
      gj_timerDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_sample_start_
      -- 
    timerDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(9) & timerDaemon_CP_9188_elements(12);
      gj_timerDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	38 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_update_start_
      -- 
    timerDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(9) & timerDaemon_CP_9188_elements(38);
      gj_timerDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_sample_completed__ps
      -- 
    -- Element group timerDaemon_CP_9188_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	37 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_update_completed__ps
      -- 
    -- Element group timerDaemon_CP_9188_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_loopback_trigger
      -- 
    timerDaemon_CP_9188_elements(19) <= timerDaemon_CP_9188_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_loopback_sample_req_ps
      -- 
    phi_stmt_4046_loopback_sample_req_9227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4046_loopback_sample_req_9227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(20), ack => phi_stmt_4046_req_0); -- 
    -- Element group timerDaemon_CP_9188_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_entry_trigger
      -- 
    timerDaemon_CP_9188_elements(21) <= timerDaemon_CP_9188_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_entry_sample_req_ps
      -- 
    phi_stmt_4046_entry_sample_req_9230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_4046_entry_sample_req_9230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(22), ack => phi_stmt_4046_req_1); -- 
    -- Element group timerDaemon_CP_9188_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4046_phi_mux_ack_ps
      -- 
    phi_stmt_4046_phi_mux_ack_9233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_4046_ack_0, ack => timerDaemon_CP_9188_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Sample/req
      -- 
    req_9246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(24), ack => nCOUNTER_4059_4048_buf_req_0); -- 
    -- Element group timerDaemon_CP_9188_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_update_start_
      -- CP-element group 25: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Update/req
      -- 
    req_9251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(25), ack => nCOUNTER_4059_4048_buf_req_1); -- 
    -- Element group timerDaemon_CP_9188_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Sample/ack
      -- 
    ack_9247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_4059_4048_buf_ack_0, ack => timerDaemon_CP_9188_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/R_nCOUNTER_4048_Update/ack
      -- 
    ack_9252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_4059_4048_buf_ack_1, ack => timerDaemon_CP_9188_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_sample_completed_
      -- 
    -- Element group timerDaemon_CP_9188_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_update_start_
      -- 
    -- Element group timerDaemon_CP_9188_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_update_completed__ps
      -- 
    timerDaemon_CP_9188_elements(30) <= timerDaemon_CP_9188_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/type_cast_4050_update_completed_
      -- 
    -- Element group timerDaemon_CP_9188_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => timerDaemon_CP_9188_elements(29), ack => timerDaemon_CP_9188_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	9 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	38 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	13 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4051_update_start_
      -- 
    timerDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(9) & timerDaemon_CP_9188_elements(38);
      gj_timerDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	11 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Sample/rr
      -- 
    rr_9273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_9273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(33), ack => RPIPE_timer_req_4053_inst_req_0); -- 
    timerDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(11) & timerDaemon_CP_9188_elements(36);
      gj_timerDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: 	13 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_update_start_
      -- CP-element group 34: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Update/cr
      -- 
    cr_9278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_9278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(34), ack => RPIPE_timer_req_4053_inst_req_1); -- 
    timerDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(35) & timerDaemon_CP_9188_elements(13);
      gj_timerDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: 	12 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Sample/ra
      -- 
    ra_9274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_4053_inst_ack_0, ack => timerDaemon_CP_9188_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: 	14 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/phi_stmt_4051_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/RPIPE_timer_req_4053_Update/ca
      -- 
    ca_9279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_timer_req_4053_inst_ack_1, ack => timerDaemon_CP_9188_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	18 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Sample/req
      -- CP-element group 37: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Sample/$entry
      -- 
    req_9287_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9287_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(37), ack => WPIPE_timer_resp_4061_inst_req_0); -- 
    timerDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(36) & timerDaemon_CP_9188_elements(18) & timerDaemon_CP_9188_elements(39);
      gj_timerDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	32 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Sample/ack
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Update/req
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_update_start_
      -- 
    ack_9288_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_4061_inst_ack_0, ack => timerDaemon_CP_9188_elements(38)); -- 
    req_9292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_9292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => timerDaemon_CP_9188_elements(38), ack => WPIPE_timer_resp_4061_inst_req_1); -- 
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/WPIPE_timer_resp_4061_update_completed_
      -- 
    ack_9293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_timer_resp_4061_inst_ack_1, ack => timerDaemon_CP_9188_elements(39)); -- 
    -- CP-element group 40:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	10 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group timerDaemon_CP_9188_elements(40) is a control-delay.
    cp_element_40_delay: control_delay_element  generic map(name => " 40_delay", delay_value => 1)  port map(req => timerDaemon_CP_9188_elements(9), ack => timerDaemon_CP_9188_elements(40), clk => clk, reset =>reset);
    -- CP-element group 41:  join  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: 	12 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	6 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_4043/do_while_stmt_4044/do_while_stmt_4044_loop_body/$exit
      -- 
    timerDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "timerDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= timerDaemon_CP_9188_elements(39) & timerDaemon_CP_9188_elements(12);
      gj_timerDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => timerDaemon_CP_9188_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	5 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_exit/$exit
      -- CP-element group 42: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_exit/ack
      -- 
    ack_9298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_4044_branch_ack_0, ack => timerDaemon_CP_9188_elements(42)); -- 
    -- CP-element group 43:  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	5 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_taken/$exit
      -- CP-element group 43: 	 branch_block_stmt_4043/do_while_stmt_4044/loop_taken/ack
      -- 
    ack_9302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_4044_branch_ack_1, ack => timerDaemon_CP_9188_elements(43)); -- 
    -- CP-element group 44:  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	3 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	1 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_4043/do_while_stmt_4044/$exit
      -- 
    timerDaemon_CP_9188_elements(44) <= timerDaemon_CP_9188_elements(3);
    timerDaemon_do_while_stmt_4044_terminator_9303: loop_terminator -- 
      generic map (name => " timerDaemon_do_while_stmt_4044_terminator_9303", max_iterations_in_flight =>7) 
      port map(loop_body_exit => timerDaemon_CP_9188_elements(6),loop_continue => timerDaemon_CP_9188_elements(43),loop_terminate => timerDaemon_CP_9188_elements(42),loop_back => timerDaemon_CP_9188_elements(4),loop_exit => timerDaemon_CP_9188_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_4046_phi_seq_9261_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= timerDaemon_CP_9188_elements(19);
      timerDaemon_CP_9188_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= timerDaemon_CP_9188_elements(26);
      timerDaemon_CP_9188_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= timerDaemon_CP_9188_elements(27);
      timerDaemon_CP_9188_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= timerDaemon_CP_9188_elements(21);
      timerDaemon_CP_9188_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= timerDaemon_CP_9188_elements(28);
      timerDaemon_CP_9188_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= timerDaemon_CP_9188_elements(30);
      timerDaemon_CP_9188_elements(22) <= phi_mux_reqs(1);
      phi_stmt_4046_phi_seq_9261 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_4046_phi_seq_9261") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => timerDaemon_CP_9188_elements(11), 
          phi_sample_ack => timerDaemon_CP_9188_elements(17), 
          phi_update_req => timerDaemon_CP_9188_elements(13), 
          phi_update_ack => timerDaemon_CP_9188_elements(18), 
          phi_mux_ack => timerDaemon_CP_9188_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_9213_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= timerDaemon_CP_9188_elements(7);
        preds(1)  <= timerDaemon_CP_9188_elements(8);
        entry_tmerge_9213 : transition_merge -- 
          generic map(name => " entry_tmerge_9213")
          port map (preds => preds, symbol_out => timerDaemon_CP_9188_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal COUNTER_4046 : std_logic_vector(63 downto 0);
    signal RPIPE_timer_req_4053_wire : std_logic_vector(0 downto 0);
    signal konst_4057_wire_constant : std_logic_vector(63 downto 0);
    signal konst_4065_wire_constant : std_logic_vector(0 downto 0);
    signal nCOUNTER_4059 : std_logic_vector(63 downto 0);
    signal nCOUNTER_4059_4048_buffered : std_logic_vector(63 downto 0);
    signal req_4051 : std_logic_vector(0 downto 0);
    signal type_cast_4050_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_4057_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    konst_4065_wire_constant <= "1";
    type_cast_4050_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_4046: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nCOUNTER_4059_4048_buffered & type_cast_4050_wire_constant;
      req <= phi_stmt_4046_req_0 & phi_stmt_4046_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_4046",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_4046_ack_0,
          idata => idata,
          odata => COUNTER_4046,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_4046
    nCOUNTER_4059_4048_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_4059_4048_buf_req_0;
      nCOUNTER_4059_4048_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_4059_4048_buf_req_1;
      nCOUNTER_4059_4048_buf_ack_1<= rack(0);
      nCOUNTER_4059_4048_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_4059_4048_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_4059,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_4059_4048_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_4051
    process(RPIPE_timer_req_4053_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := RPIPE_timer_req_4053_wire(0 downto 0);
      req_4051 <= tmp_var; -- 
    end process;
    do_while_stmt_4044_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_4065_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_4044_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_4044_branch_req_0,
          ack0 => do_while_stmt_4044_branch_ack_0,
          ack1 => do_while_stmt_4044_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u64_u64_4058_inst
    process(COUNTER_4046) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_4046, konst_4057_wire_constant, tmp_var);
      nCOUNTER_4059 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_timer_req_4053_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_timer_req_4053_inst_req_0;
      RPIPE_timer_req_4053_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_timer_req_4053_inst_req_1;
      RPIPE_timer_req_4053_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_timer_req_4053_wire <= data_out(0 downto 0);
      timer_req_read_0_gI: SplitGuardInterface generic map(name => "timer_req_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      timer_req_read_0: InputPortRevised -- 
        generic map ( name => "timer_req_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => timer_req_pipe_read_req(0),
          oack => timer_req_pipe_read_ack(0),
          odata => timer_req_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_timer_resp_4061_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_timer_resp_4061_inst_req_0;
      WPIPE_timer_resp_4061_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_timer_resp_4061_inst_req_1;
      WPIPE_timer_resp_4061_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= req_4051(0);
      data_in <= COUNTER_4046;
      timer_resp_write_0_gI: SplitGuardInterface generic map(name => "timer_resp_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      timer_resp_write_0: OutputPortRevised -- 
        generic map ( name => "timer_resp", data_width => 64, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => timer_resp_pipe_write_req(0),
          oack => timer_resp_pipe_write_ack(0),
          odata => timer_resp_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end timerDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    maxpool_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    maxpool_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    maxpool_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    maxpool_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    maxpool_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(27 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(37 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(127 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(2 downto 0);
  -- declarations related to module access_T
  component access_T is -- 
    generic (tag_length : integer); 
    port ( -- 
      row_in : in  std_logic_vector(15 downto 0);
      chl_in : in  std_logic_vector(15 downto 0);
      ct : in  std_logic_vector(15 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      input_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
      input_pipe4_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module access_T
  signal access_T_row_in :  std_logic_vector(15 downto 0);
  signal access_T_chl_in :  std_logic_vector(15 downto 0);
  signal access_T_ct :  std_logic_vector(15 downto 0);
  signal access_T_in_args    : std_logic_vector(47 downto 0);
  signal access_T_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal access_T_tag_out   : std_logic_vector(1 downto 0);
  signal access_T_start_req : std_logic;
  signal access_T_start_ack : std_logic;
  signal access_T_fin_req   : std_logic;
  signal access_T_fin_ack : std_logic;
  -- caller side aggregated signals for module access_T
  signal access_T_call_reqs: std_logic_vector(0 downto 0);
  signal access_T_call_acks: std_logic_vector(0 downto 0);
  signal access_T_return_reqs: std_logic_vector(0 downto 0);
  signal access_T_return_acks: std_logic_vector(0 downto 0);
  signal access_T_call_data: std_logic_vector(47 downto 0);
  signal access_T_call_tag: std_logic_vector(0 downto 0);
  signal access_T_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module convolution3D
  component convolution3D is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      maxpool_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      num_out_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      timer_call_reqs : out  std_logic_vector(0 downto 0);
      timer_call_acks : in   std_logic_vector(0 downto 0);
      timer_call_tag  :  out  std_logic_vector(1 downto 0);
      timer_return_reqs : out  std_logic_vector(0 downto 0);
      timer_return_acks : in   std_logic_vector(0 downto 0);
      timer_return_data : in   std_logic_vector(63 downto 0);
      timer_return_tag :  in   std_logic_vector(1 downto 0);
      access_T_call_reqs : out  std_logic_vector(0 downto 0);
      access_T_call_acks : in   std_logic_vector(0 downto 0);
      access_T_call_data : out  std_logic_vector(47 downto 0);
      access_T_call_tag  :  out  std_logic_vector(0 downto 0);
      access_T_return_reqs : out  std_logic_vector(0 downto 0);
      access_T_return_acks : in   std_logic_vector(0 downto 0);
      access_T_return_tag :  in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_call_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_call_data : out  std_logic_vector(47 downto 0);
      loadKernelChannel_call_tag  :  out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_reqs : out  std_logic_vector(0 downto 0);
      loadKernelChannel_return_acks : in   std_logic_vector(0 downto 0);
      loadKernelChannel_return_tag :  in   std_logic_vector(0 downto 0);
      sendB_call_reqs : out  std_logic_vector(0 downto 0);
      sendB_call_acks : in   std_logic_vector(0 downto 0);
      sendB_call_data : out  std_logic_vector(31 downto 0);
      sendB_call_tag  :  out  std_logic_vector(0 downto 0);
      sendB_return_reqs : out  std_logic_vector(0 downto 0);
      sendB_return_acks : in   std_logic_vector(0 downto 0);
      sendB_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolution3D
  signal convolution3D_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolution3D_tag_out   : std_logic_vector(1 downto 0);
  signal convolution3D_start_req : std_logic;
  signal convolution3D_start_ack : std_logic;
  signal convolution3D_fin_req   : std_logic;
  signal convolution3D_fin_ack : std_logic;
  -- declarations related to module convolve
  component convolve is -- 
    generic (tag_length : integer); 
    port ( -- 
      input_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe2_pipe_read_data : in   std_logic_vector(63 downto 0);
      input_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe3_pipe_read_data : in   std_logic_vector(63 downto 0);
      input_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe1_pipe_read_data : in   std_logic_vector(63 downto 0);
      kernel_pipe2_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_read_data : in   std_logic_vector(63 downto 0);
      kernel_pipe3_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_read_data : in   std_logic_vector(63 downto 0);
      input_pipe4_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_pipe4_pipe_read_data : in   std_logic_vector(63 downto 0);
      kernel_pipe1_pipe_read_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_read_data : in   std_logic_vector(63 downto 0);
      num_out_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      num_out_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      size_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_read_data : in   std_logic_vector(15 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      output_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convolve
  signal convolve_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convolve_tag_out   : std_logic_vector(1 downto 0);
  signal convolve_start_req : std_logic;
  signal convolve_start_ack : std_logic;
  signal convolve_fin_req   : std_logic;
  signal convolve_fin_ack : std_logic;
  -- declarations related to module loadKernelChannel
  component loadKernelChannel is -- 
    generic (tag_length : integer); 
    port ( -- 
      start_add : in  std_logic_vector(31 downto 0);
      num_chl : in  std_logic_vector(15 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(1 downto 0);
      input_done_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      kernel_pipe2_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe2_pipe_write_data : out  std_logic_vector(63 downto 0);
      kernel_pipe3_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe3_pipe_write_data : out  std_logic_vector(63 downto 0);
      kernel_pipe1_pipe_write_req : out  std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_ack : in   std_logic_vector(0 downto 0);
      kernel_pipe1_pipe_write_data : out  std_logic_vector(63 downto 0);
      size_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      size_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      size_pipe_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadKernelChannel
  signal loadKernelChannel_start_add :  std_logic_vector(31 downto 0);
  signal loadKernelChannel_num_chl :  std_logic_vector(15 downto 0);
  signal loadKernelChannel_in_args    : std_logic_vector(47 downto 0);
  signal loadKernelChannel_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadKernelChannel_tag_out   : std_logic_vector(1 downto 0);
  signal loadKernelChannel_start_req : std_logic;
  signal loadKernelChannel_start_ack : std_logic;
  signal loadKernelChannel_fin_req   : std_logic;
  signal loadKernelChannel_fin_ack : std_logic;
  -- caller side aggregated signals for module loadKernelChannel
  signal loadKernelChannel_call_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_reqs: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_acks: std_logic_vector(0 downto 0);
  signal loadKernelChannel_call_data: std_logic_vector(47 downto 0);
  signal loadKernelChannel_call_tag: std_logic_vector(0 downto 0);
  signal loadKernelChannel_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendB
  component sendB is -- 
    generic (tag_length : integer); 
    port ( -- 
      size : in  std_logic_vector(31 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      maxpool_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      maxpool_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendB
  signal sendB_size :  std_logic_vector(31 downto 0);
  signal sendB_in_args    : std_logic_vector(31 downto 0);
  signal sendB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendB_tag_out   : std_logic_vector(1 downto 0);
  signal sendB_start_req : std_logic;
  signal sendB_start_ack : std_logic;
  signal sendB_fin_req   : std_logic;
  signal sendB_fin_ack : std_logic;
  -- caller side aggregated signals for module sendB
  signal sendB_call_reqs: std_logic_vector(0 downto 0);
  signal sendB_call_acks: std_logic_vector(0 downto 0);
  signal sendB_return_reqs: std_logic_vector(0 downto 0);
  signal sendB_return_acks: std_logic_vector(0 downto 0);
  signal sendB_call_data: std_logic_vector(31 downto 0);
  signal sendB_call_tag: std_logic_vector(0 downto 0);
  signal sendB_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendModule
  component sendModule is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_req : out  std_logic_vector(1 downto 0);
      output_pipe_pipe_read_ack : in   std_logic_vector(1 downto 0);
      output_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      input_done_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      input_done_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendModule
  signal sendModule_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendModule_tag_out   : std_logic_vector(1 downto 0);
  signal sendModule_start_req : std_logic;
  signal sendModule_start_ack : std_logic;
  signal sendModule_fin_req   : std_logic;
  signal sendModule_fin_ack : std_logic;
  -- declarations related to module timer
  component timer is -- 
    generic (tag_length : integer); 
    port ( -- 
      T : out  std_logic_vector(63 downto 0);
      timer_resp_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_read_data : in   std_logic_vector(63 downto 0);
      timer_req_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_write_data : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timer
  signal timer_T :  std_logic_vector(63 downto 0);
  signal timer_out_args   : std_logic_vector(63 downto 0);
  signal timer_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal timer_tag_out   : std_logic_vector(2 downto 0);
  signal timer_start_req : std_logic;
  signal timer_start_ack : std_logic;
  signal timer_fin_req   : std_logic;
  signal timer_fin_ack : std_logic;
  -- caller side aggregated signals for module timer
  signal timer_call_reqs: std_logic_vector(0 downto 0);
  signal timer_call_acks: std_logic_vector(0 downto 0);
  signal timer_return_reqs: std_logic_vector(0 downto 0);
  signal timer_return_acks: std_logic_vector(0 downto 0);
  signal timer_call_tag: std_logic_vector(1 downto 0);
  signal timer_return_data: std_logic_vector(63 downto 0);
  signal timer_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module timerDaemon
  component timerDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      timer_req_pipe_read_req : out  std_logic_vector(0 downto 0);
      timer_req_pipe_read_ack : in   std_logic_vector(0 downto 0);
      timer_req_pipe_read_data : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_req : out  std_logic_vector(0 downto 0);
      timer_resp_pipe_write_ack : in   std_logic_vector(0 downto 0);
      timer_resp_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module timerDaemon
  signal timerDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal timerDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal timerDaemon_start_req : std_logic;
  signal timerDaemon_start_ack : std_logic;
  signal timerDaemon_fin_req   : std_logic;
  signal timerDaemon_fin_ack : std_logic;
  -- aggregate signals for write to pipe input_done_pipe
  signal input_done_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe input_done_pipe
  signal input_done_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal input_done_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal input_done_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe input_pipe1
  signal input_pipe1_pipe_write_data: std_logic_vector(63 downto 0);
  signal input_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe1
  signal input_pipe1_pipe_read_data: std_logic_vector(63 downto 0);
  signal input_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe2
  signal input_pipe2_pipe_write_data: std_logic_vector(63 downto 0);
  signal input_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe2
  signal input_pipe2_pipe_read_data: std_logic_vector(63 downto 0);
  signal input_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe3
  signal input_pipe3_pipe_write_data: std_logic_vector(63 downto 0);
  signal input_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe3
  signal input_pipe3_pipe_read_data: std_logic_vector(63 downto 0);
  signal input_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe input_pipe4
  signal input_pipe4_pipe_write_data: std_logic_vector(63 downto 0);
  signal input_pipe4_pipe_write_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe input_pipe4
  signal input_pipe4_pipe_read_data: std_logic_vector(63 downto 0);
  signal input_pipe4_pipe_read_req: std_logic_vector(0 downto 0);
  signal input_pipe4_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe1
  signal kernel_pipe1_pipe_write_data: std_logic_vector(63 downto 0);
  signal kernel_pipe1_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe1
  signal kernel_pipe1_pipe_read_data: std_logic_vector(63 downto 0);
  signal kernel_pipe1_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe1_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe2
  signal kernel_pipe2_pipe_write_data: std_logic_vector(63 downto 0);
  signal kernel_pipe2_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe2
  signal kernel_pipe2_pipe_read_data: std_logic_vector(63 downto 0);
  signal kernel_pipe2_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe2_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe kernel_pipe3
  signal kernel_pipe3_pipe_write_data: std_logic_vector(63 downto 0);
  signal kernel_pipe3_pipe_write_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe kernel_pipe3
  signal kernel_pipe3_pipe_read_data: std_logic_vector(63 downto 0);
  signal kernel_pipe3_pipe_read_req: std_logic_vector(0 downto 0);
  signal kernel_pipe3_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe maxpool_input_pipe
  signal maxpool_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal maxpool_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal maxpool_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe maxpool_output_pipe
  signal maxpool_output_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal maxpool_output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal maxpool_output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe num_out_pipe
  signal num_out_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe num_out_pipe
  signal num_out_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal num_out_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal num_out_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe output_pipe
  signal output_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe output_pipe
  signal output_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal output_pipe_pipe_read_req: std_logic_vector(1 downto 0);
  signal output_pipe_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe size_pipe
  signal size_pipe_pipe_write_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe size_pipe
  signal size_pipe_pipe_read_data: std_logic_vector(15 downto 0);
  signal size_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal size_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_req
  signal timer_req_pipe_write_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_req
  signal timer_req_pipe_read_data: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_req_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe timer_resp
  signal timer_resp_pipe_write_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_write_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe timer_resp
  signal timer_resp_pipe_read_data: std_logic_vector(63 downto 0);
  signal timer_resp_pipe_read_req: std_logic_vector(0 downto 0);
  signal timer_resp_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module access_T
  access_T_row_in <= access_T_in_args(47 downto 32);
  access_T_chl_in <= access_T_in_args(31 downto 16);
  access_T_ct <= access_T_in_args(15 downto 0);
  -- call arbiter for module access_T
  access_T_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => access_T_call_reqs,
      call_acks => access_T_call_acks,
      return_reqs => access_T_return_reqs,
      return_acks => access_T_return_acks,
      call_data  => access_T_call_data,
      call_tag  => access_T_call_tag,
      return_tag  => access_T_return_tag,
      call_mtag => access_T_tag_in,
      return_mtag => access_T_tag_out,
      call_mreq => access_T_start_req,
      call_mack => access_T_start_ack,
      return_mreq => access_T_fin_req,
      return_mack => access_T_fin_ack,
      call_mdata => access_T_in_args,
      clk => clk, 
      reset => reset --
    ); --
  access_T_instance:access_T-- 
    generic map(tag_length => 2)
    port map(-- 
      row_in => access_T_row_in,
      chl_in => access_T_chl_in,
      ct => access_T_ct,
      start_req => access_T_start_req,
      start_ack => access_T_start_ack,
      fin_req => access_T_fin_req,
      fin_ack => access_T_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      input_pipe2_pipe_write_req => input_pipe2_pipe_write_req(0 downto 0),
      input_pipe2_pipe_write_ack => input_pipe2_pipe_write_ack(0 downto 0),
      input_pipe2_pipe_write_data => input_pipe2_pipe_write_data(63 downto 0),
      input_pipe3_pipe_write_req => input_pipe3_pipe_write_req(0 downto 0),
      input_pipe3_pipe_write_ack => input_pipe3_pipe_write_ack(0 downto 0),
      input_pipe3_pipe_write_data => input_pipe3_pipe_write_data(63 downto 0),
      input_pipe1_pipe_write_req => input_pipe1_pipe_write_req(0 downto 0),
      input_pipe1_pipe_write_ack => input_pipe1_pipe_write_ack(0 downto 0),
      input_pipe1_pipe_write_data => input_pipe1_pipe_write_data(63 downto 0),
      input_pipe4_pipe_write_req => input_pipe4_pipe_write_req(0 downto 0),
      input_pipe4_pipe_write_ack => input_pipe4_pipe_write_ack(0 downto 0),
      input_pipe4_pipe_write_data => input_pipe4_pipe_write_data(63 downto 0),
      tag_in => access_T_tag_in,
      tag_out => access_T_tag_out-- 
    ); -- 
  -- module convolution3D
  convolution3D_instance:convolution3D-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolution3D_start_req,
      start_ack => convolution3D_start_ack,
      fin_req => convolution3D_fin_req,
      fin_ack => convolution3D_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(13 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(63 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(18 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(13 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(0 downto 0),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(0 downto 0),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(7 downto 0),
      maxpool_input_pipe_pipe_read_req => maxpool_input_pipe_pipe_read_req(0 downto 0),
      maxpool_input_pipe_pipe_read_ack => maxpool_input_pipe_pipe_read_ack(0 downto 0),
      maxpool_input_pipe_pipe_read_data => maxpool_input_pipe_pipe_read_data(7 downto 0),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(0 downto 0),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(0 downto 0),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(7 downto 0),
      num_out_pipe_pipe_write_req => num_out_pipe_pipe_write_req(0 downto 0),
      num_out_pipe_pipe_write_ack => num_out_pipe_pipe_write_ack(0 downto 0),
      num_out_pipe_pipe_write_data => num_out_pipe_pipe_write_data(15 downto 0),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(1 downto 1),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(1 downto 1),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(31 downto 16),
      access_T_call_reqs => access_T_call_reqs(0 downto 0),
      access_T_call_acks => access_T_call_acks(0 downto 0),
      access_T_call_data => access_T_call_data(47 downto 0),
      access_T_call_tag => access_T_call_tag(0 downto 0),
      access_T_return_reqs => access_T_return_reqs(0 downto 0),
      access_T_return_acks => access_T_return_acks(0 downto 0),
      access_T_return_tag => access_T_return_tag(0 downto 0),
      timer_call_reqs => timer_call_reqs(0 downto 0),
      timer_call_acks => timer_call_acks(0 downto 0),
      timer_call_tag => timer_call_tag(1 downto 0),
      timer_return_reqs => timer_return_reqs(0 downto 0),
      timer_return_acks => timer_return_acks(0 downto 0),
      timer_return_data => timer_return_data(63 downto 0),
      timer_return_tag => timer_return_tag(1 downto 0),
      loadKernelChannel_call_reqs => loadKernelChannel_call_reqs(0 downto 0),
      loadKernelChannel_call_acks => loadKernelChannel_call_acks(0 downto 0),
      loadKernelChannel_call_data => loadKernelChannel_call_data(47 downto 0),
      loadKernelChannel_call_tag => loadKernelChannel_call_tag(0 downto 0),
      loadKernelChannel_return_reqs => loadKernelChannel_return_reqs(0 downto 0),
      loadKernelChannel_return_acks => loadKernelChannel_return_acks(0 downto 0),
      loadKernelChannel_return_tag => loadKernelChannel_return_tag(0 downto 0),
      sendB_call_reqs => sendB_call_reqs(0 downto 0),
      sendB_call_acks => sendB_call_acks(0 downto 0),
      sendB_call_data => sendB_call_data(31 downto 0),
      sendB_call_tag => sendB_call_tag(0 downto 0),
      sendB_return_reqs => sendB_return_reqs(0 downto 0),
      sendB_return_acks => sendB_return_acks(0 downto 0),
      sendB_return_tag => sendB_return_tag(0 downto 0),
      tag_in => convolution3D_tag_in,
      tag_out => convolution3D_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolution3D_tag_in <= (others => '0');
  convolution3D_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolution3D_start_req, start_ack => convolution3D_start_ack,  fin_req => convolution3D_fin_req,  fin_ack => convolution3D_fin_ack);
  -- module convolve
  convolve_instance:convolve-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convolve_start_req,
      start_ack => convolve_start_ack,
      fin_req => convolve_fin_req,
      fin_ack => convolve_fin_ack,
      clk => clk,
      reset => reset,
      input_pipe2_pipe_read_req => input_pipe2_pipe_read_req(0 downto 0),
      input_pipe2_pipe_read_ack => input_pipe2_pipe_read_ack(0 downto 0),
      input_pipe2_pipe_read_data => input_pipe2_pipe_read_data(63 downto 0),
      input_pipe3_pipe_read_req => input_pipe3_pipe_read_req(0 downto 0),
      input_pipe3_pipe_read_ack => input_pipe3_pipe_read_ack(0 downto 0),
      input_pipe3_pipe_read_data => input_pipe3_pipe_read_data(63 downto 0),
      input_pipe1_pipe_read_req => input_pipe1_pipe_read_req(0 downto 0),
      input_pipe1_pipe_read_ack => input_pipe1_pipe_read_ack(0 downto 0),
      input_pipe1_pipe_read_data => input_pipe1_pipe_read_data(63 downto 0),
      kernel_pipe2_pipe_read_req => kernel_pipe2_pipe_read_req(0 downto 0),
      kernel_pipe2_pipe_read_ack => kernel_pipe2_pipe_read_ack(0 downto 0),
      kernel_pipe2_pipe_read_data => kernel_pipe2_pipe_read_data(63 downto 0),
      kernel_pipe3_pipe_read_req => kernel_pipe3_pipe_read_req(0 downto 0),
      kernel_pipe3_pipe_read_ack => kernel_pipe3_pipe_read_ack(0 downto 0),
      kernel_pipe3_pipe_read_data => kernel_pipe3_pipe_read_data(63 downto 0),
      input_pipe4_pipe_read_req => input_pipe4_pipe_read_req(0 downto 0),
      input_pipe4_pipe_read_ack => input_pipe4_pipe_read_ack(0 downto 0),
      input_pipe4_pipe_read_data => input_pipe4_pipe_read_data(63 downto 0),
      kernel_pipe1_pipe_read_req => kernel_pipe1_pipe_read_req(0 downto 0),
      kernel_pipe1_pipe_read_ack => kernel_pipe1_pipe_read_ack(0 downto 0),
      kernel_pipe1_pipe_read_data => kernel_pipe1_pipe_read_data(63 downto 0),
      num_out_pipe_pipe_read_req => num_out_pipe_pipe_read_req(0 downto 0),
      num_out_pipe_pipe_read_ack => num_out_pipe_pipe_read_ack(0 downto 0),
      num_out_pipe_pipe_read_data => num_out_pipe_pipe_read_data(15 downto 0),
      size_pipe_pipe_read_req => size_pipe_pipe_read_req(0 downto 0),
      size_pipe_pipe_read_ack => size_pipe_pipe_read_ack(0 downto 0),
      size_pipe_pipe_read_data => size_pipe_pipe_read_data(15 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(1 downto 1),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(1 downto 1),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(15 downto 8),
      output_pipe_pipe_write_req => output_pipe_pipe_write_req(0 downto 0),
      output_pipe_pipe_write_ack => output_pipe_pipe_write_ack(0 downto 0),
      output_pipe_pipe_write_data => output_pipe_pipe_write_data(15 downto 0),
      tag_in => convolve_tag_in,
      tag_out => convolve_tag_out-- 
    ); -- 
  -- module will be run forever 
  convolve_tag_in <= (others => '0');
  convolve_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convolve_start_req, start_ack => convolve_start_ack,  fin_req => convolve_fin_req,  fin_ack => convolve_fin_ack);
  -- module loadKernelChannel
  loadKernelChannel_start_add <= loadKernelChannel_in_args(47 downto 16);
  loadKernelChannel_num_chl <= loadKernelChannel_in_args(15 downto 0);
  -- call arbiter for module loadKernelChannel
  loadKernelChannel_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 48,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadKernelChannel_call_reqs,
      call_acks => loadKernelChannel_call_acks,
      return_reqs => loadKernelChannel_return_reqs,
      return_acks => loadKernelChannel_return_acks,
      call_data  => loadKernelChannel_call_data,
      call_tag  => loadKernelChannel_call_tag,
      return_tag  => loadKernelChannel_return_tag,
      call_mtag => loadKernelChannel_tag_in,
      return_mtag => loadKernelChannel_tag_out,
      call_mreq => loadKernelChannel_start_req,
      call_mack => loadKernelChannel_start_ack,
      return_mreq => loadKernelChannel_fin_req,
      return_mack => loadKernelChannel_fin_ack,
      call_mdata => loadKernelChannel_in_args,
      clk => clk, 
      reset => reset --
    ); --
  loadKernelChannel_instance:loadKernelChannel-- 
    generic map(tag_length => 2)
    port map(-- 
      start_add => loadKernelChannel_start_add,
      num_chl => loadKernelChannel_num_chl,
      start_req => loadKernelChannel_start_req,
      start_ack => loadKernelChannel_start_ack,
      fin_req => loadKernelChannel_fin_req,
      fin_ack => loadKernelChannel_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(18 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(1 downto 0),
      input_done_pipe_pipe_read_req => input_done_pipe_pipe_read_req(1 downto 1),
      input_done_pipe_pipe_read_ack => input_done_pipe_pipe_read_ack(1 downto 1),
      input_done_pipe_pipe_read_data => input_done_pipe_pipe_read_data(15 downto 8),
      kernel_pipe2_pipe_write_req => kernel_pipe2_pipe_write_req(0 downto 0),
      kernel_pipe2_pipe_write_ack => kernel_pipe2_pipe_write_ack(0 downto 0),
      kernel_pipe2_pipe_write_data => kernel_pipe2_pipe_write_data(63 downto 0),
      kernel_pipe3_pipe_write_req => kernel_pipe3_pipe_write_req(0 downto 0),
      kernel_pipe3_pipe_write_ack => kernel_pipe3_pipe_write_ack(0 downto 0),
      kernel_pipe3_pipe_write_data => kernel_pipe3_pipe_write_data(63 downto 0),
      kernel_pipe1_pipe_write_req => kernel_pipe1_pipe_write_req(0 downto 0),
      kernel_pipe1_pipe_write_ack => kernel_pipe1_pipe_write_ack(0 downto 0),
      kernel_pipe1_pipe_write_data => kernel_pipe1_pipe_write_data(63 downto 0),
      size_pipe_pipe_write_req => size_pipe_pipe_write_req(0 downto 0),
      size_pipe_pipe_write_ack => size_pipe_pipe_write_ack(0 downto 0),
      size_pipe_pipe_write_data => size_pipe_pipe_write_data(15 downto 0),
      tag_in => loadKernelChannel_tag_in,
      tag_out => loadKernelChannel_tag_out-- 
    ); -- 
  -- module sendB
  sendB_size <= sendB_in_args(31 downto 0);
  -- call arbiter for module sendB
  sendB_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendB_call_reqs,
      call_acks => sendB_call_acks,
      return_reqs => sendB_return_reqs,
      return_acks => sendB_return_acks,
      call_data  => sendB_call_data,
      call_tag  => sendB_call_tag,
      return_tag  => sendB_return_tag,
      call_mtag => sendB_tag_in,
      return_mtag => sendB_tag_out,
      call_mreq => sendB_start_req,
      call_mack => sendB_start_ack,
      return_mreq => sendB_fin_req,
      return_mack => sendB_fin_ack,
      call_mdata => sendB_in_args,
      clk => clk, 
      reset => reset --
    ); --
  sendB_instance:sendB-- 
    generic map(tag_length => 2)
    port map(-- 
      size => sendB_size,
      start_req => sendB_start_req,
      start_ack => sendB_start_ack,
      fin_req => sendB_fin_req,
      fin_ack => sendB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(37 downto 19),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 2),
      maxpool_output_pipe_pipe_write_req => maxpool_output_pipe_pipe_write_req(1 downto 1),
      maxpool_output_pipe_pipe_write_ack => maxpool_output_pipe_pipe_write_ack(1 downto 1),
      maxpool_output_pipe_pipe_write_data => maxpool_output_pipe_pipe_write_data(15 downto 8),
      tag_in => sendB_tag_in,
      tag_out => sendB_tag_out-- 
    ); -- 
  -- module sendModule
  sendModule_instance:sendModule-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendModule_start_req,
      start_ack => sendModule_start_ack,
      fin_req => sendModule_fin_req,
      fin_ack => sendModule_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(18 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(1 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(13 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(63 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(18 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(1 downto 0),
      output_pipe_pipe_read_req => output_pipe_pipe_read_req(1 downto 0),
      output_pipe_pipe_read_ack => output_pipe_pipe_read_ack(1 downto 0),
      output_pipe_pipe_read_data => output_pipe_pipe_read_data(31 downto 0),
      input_done_pipe_pipe_write_req => input_done_pipe_pipe_write_req(0 downto 0),
      input_done_pipe_pipe_write_ack => input_done_pipe_pipe_write_ack(0 downto 0),
      input_done_pipe_pipe_write_data => input_done_pipe_pipe_write_data(7 downto 0),
      tag_in => sendModule_tag_in,
      tag_out => sendModule_tag_out-- 
    ); -- 
  -- module will be run forever 
  sendModule_tag_in <= (others => '0');
  sendModule_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => sendModule_start_req, start_ack => sendModule_start_ack,  fin_req => sendModule_fin_req,  fin_ack => sendModule_fin_ack);
  -- module timer
  timer_out_args <= timer_T ;
  -- call arbiter for module timer
  timer_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => timer_call_reqs,
      call_acks => timer_call_acks,
      return_reqs => timer_return_reqs,
      return_acks => timer_return_acks,
      call_tag  => timer_call_tag,
      return_tag  => timer_return_tag,
      call_mtag => timer_tag_in,
      return_mtag => timer_tag_out,
      return_data =>timer_return_data,
      call_mreq => timer_start_req,
      call_mack => timer_start_ack,
      return_mreq => timer_fin_req,
      return_mack => timer_fin_ack,
      return_mdata => timer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  timer_instance:timer-- 
    generic map(tag_length => 3)
    port map(-- 
      T => timer_T,
      start_req => timer_start_req,
      start_ack => timer_start_ack,
      fin_req => timer_fin_req,
      fin_ack => timer_fin_ack,
      clk => clk,
      reset => reset,
      timer_resp_pipe_read_req => timer_resp_pipe_read_req(0 downto 0),
      timer_resp_pipe_read_ack => timer_resp_pipe_read_ack(0 downto 0),
      timer_resp_pipe_read_data => timer_resp_pipe_read_data(63 downto 0),
      timer_req_pipe_write_req => timer_req_pipe_write_req(0 downto 0),
      timer_req_pipe_write_ack => timer_req_pipe_write_ack(0 downto 0),
      timer_req_pipe_write_data => timer_req_pipe_write_data(0 downto 0),
      tag_in => timer_tag_in,
      tag_out => timer_tag_out-- 
    ); -- 
  -- module timerDaemon
  timerDaemon_instance:timerDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => timerDaemon_start_req,
      start_ack => timerDaemon_start_ack,
      fin_req => timerDaemon_fin_req,
      fin_ack => timerDaemon_fin_ack,
      clk => clk,
      reset => reset,
      timer_req_pipe_read_req => timer_req_pipe_read_req(0 downto 0),
      timer_req_pipe_read_ack => timer_req_pipe_read_ack(0 downto 0),
      timer_req_pipe_read_data => timer_req_pipe_read_data(0 downto 0),
      timer_resp_pipe_write_req => timer_resp_pipe_write_req(0 downto 0),
      timer_resp_pipe_write_ack => timer_resp_pipe_write_ack(0 downto 0),
      timer_resp_pipe_write_data => timer_resp_pipe_write_data(63 downto 0),
      tag_in => timerDaemon_tag_in,
      tag_out => timerDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  timerDaemon_tag_in <= (others => '0');
  timerDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => timerDaemon_start_req, start_ack => timerDaemon_start_ack,  fin_req => timerDaemon_fin_req,  fin_ack => timerDaemon_fin_ack);
  input_done_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_done_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => input_done_pipe_pipe_read_req,
      read_ack => input_done_pipe_pipe_read_ack,
      read_data => input_done_pipe_pipe_read_data,
      write_req => input_done_pipe_pipe_write_req,
      write_ack => input_done_pipe_pipe_write_ack,
      write_data => input_done_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => input_pipe1_pipe_read_req,
      read_ack => input_pipe1_pipe_read_ack,
      read_data => input_pipe1_pipe_read_data,
      write_req => input_pipe1_pipe_write_req,
      write_ack => input_pipe1_pipe_write_ack,
      write_data => input_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => input_pipe2_pipe_read_req,
      read_ack => input_pipe2_pipe_read_ack,
      read_data => input_pipe2_pipe_read_data,
      write_req => input_pipe2_pipe_write_req,
      write_ack => input_pipe2_pipe_write_ack,
      write_data => input_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => input_pipe3_pipe_read_req,
      read_ack => input_pipe3_pipe_read_ack,
      read_data => input_pipe3_pipe_read_data,
      write_req => input_pipe3_pipe_write_req,
      write_ack => input_pipe3_pipe_write_ack,
      write_data => input_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  input_pipe4_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe input_pipe4",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => input_pipe4_pipe_read_req,
      read_ack => input_pipe4_pipe_read_ack,
      read_data => input_pipe4_pipe_read_data,
      write_req => input_pipe4_pipe_write_req,
      write_ack => input_pipe4_pipe_write_ack,
      write_data => input_pipe4_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe1_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe1",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => kernel_pipe1_pipe_read_req,
      read_ack => kernel_pipe1_pipe_read_ack,
      read_data => kernel_pipe1_pipe_read_data,
      write_req => kernel_pipe1_pipe_write_req,
      write_ack => kernel_pipe1_pipe_write_ack,
      write_data => kernel_pipe1_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe2_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe2",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => kernel_pipe2_pipe_read_req,
      read_ack => kernel_pipe2_pipe_read_ack,
      read_data => kernel_pipe2_pipe_read_data,
      write_req => kernel_pipe2_pipe_write_req,
      write_ack => kernel_pipe2_pipe_write_ack,
      write_data => kernel_pipe2_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  kernel_pipe3_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe kernel_pipe3",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 64 --
    )
    port map( -- 
      read_req => kernel_pipe3_pipe_read_req,
      read_ack => kernel_pipe3_pipe_read_ack,
      read_data => kernel_pipe3_pipe_read_data,
      write_req => kernel_pipe3_pipe_write_req,
      write_ack => kernel_pipe3_pipe_write_ack,
      write_data => kernel_pipe3_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_input_pipe_pipe_read_req,
      read_ack => maxpool_input_pipe_pipe_read_ack,
      read_data => maxpool_input_pipe_pipe_read_data,
      write_req => maxpool_input_pipe_pipe_write_req,
      write_ack => maxpool_input_pipe_pipe_write_ack,
      write_data => maxpool_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  maxpool_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe maxpool_output_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => maxpool_output_pipe_pipe_read_req,
      read_ack => maxpool_output_pipe_pipe_read_ack,
      read_data => maxpool_output_pipe_pipe_read_data,
      write_req => maxpool_output_pipe_pipe_write_req,
      write_ack => maxpool_output_pipe_pipe_write_ack,
      write_data => maxpool_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  num_out_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe num_out_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => num_out_pipe_pipe_read_req,
      read_ack => num_out_pipe_pipe_read_ack,
      read_data => num_out_pipe_pipe_read_data,
      write_req => num_out_pipe_pipe_write_req,
      write_ack => num_out_pipe_pipe_write_ack,
      write_data => num_out_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe output_pipe",
      num_reads => 2,
      num_writes => 2,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 10 --
    )
    port map( -- 
      read_req => output_pipe_pipe_read_req,
      read_ack => output_pipe_pipe_read_ack,
      read_data => output_pipe_pipe_read_data,
      write_req => output_pipe_pipe_write_req,
      write_ack => output_pipe_pipe_write_ack,
      write_data => output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  size_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe size_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 4 --
    )
    port map( -- 
      read_req => size_pipe_pipe_read_req,
      read_ack => size_pipe_pipe_read_ack,
      read_data => size_pipe_pipe_read_data,
      write_req => size_pipe_pipe_write_req,
      write_ack => size_pipe_pipe_write_ack,
      write_data => size_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  timer_req_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_req",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_req_pipe_read_req,
      read_ack => timer_req_pipe_read_ack,
      read_data => timer_req_pipe_read_data,
      write_req => timer_req_pipe_write_req,
      write_ack => timer_req_pipe_write_ack,
      write_data => timer_req_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  timer_resp_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe timer_resp",
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => timer_resp_pipe_read_req,
      read_ack => timer_resp_pipe_read_ack,
      read_data => timer_resp_pipe_read_data,
      write_req => timer_resp_pipe_write_req,
      write_ack => timer_resp_pipe_write_ack,
      write_data => timer_resp_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 2,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 2,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 3,
      time_stamp_width => 17,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
