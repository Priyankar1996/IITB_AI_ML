-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTranspose is -- 
  generic (tag_length : integer); 
  port ( -- 
    Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
    testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_call_acks : in   std_logic_vector(0 downto 0);
    testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
    testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
    testConfigure_return_acks : in   std_logic_vector(0 downto 0);
    testConfigure_return_data : in   std_logic_vector(15 downto 0);
    testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
    sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_call_acks : in   std_logic_vector(0 downto 0);
    sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
    sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
    sendOutput_return_acks : in   std_logic_vector(0 downto 0);
    sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTranspose;
architecture convTranspose_arch of convTranspose is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTranspose_CP_3910_start: Boolean;
  signal convTranspose_CP_3910_symbol: Boolean;
  -- volatile/operator module components. 
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal RPIPE_Block0_done_1346_inst_req_0 : boolean;
  signal RPIPE_Block2_done_1352_inst_ack_0 : boolean;
  signal RPIPE_Block1_done_1349_inst_req_1 : boolean;
  signal RPIPE_Block1_done_1349_inst_ack_1 : boolean;
  signal WPIPE_Block0_start_1333_inst_ack_0 : boolean;
  signal RPIPE_Block3_done_1355_inst_req_0 : boolean;
  signal WPIPE_Block0_start_1333_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1355_inst_ack_0 : boolean;
  signal WPIPE_Block3_start_1342_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1336_inst_ack_1 : boolean;
  signal WPIPE_Block3_start_1342_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1352_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1346_inst_ack_0 : boolean;
  signal WPIPE_Block0_start_1333_inst_req_0 : boolean;
  signal WPIPE_Block3_start_1342_inst_ack_0 : boolean;
  signal call_stmt_1331_call_ack_1 : boolean;
  signal call_stmt_1331_call_req_1 : boolean;
  signal call_stmt_1331_call_ack_0 : boolean;
  signal WPIPE_Block3_start_1342_inst_req_0 : boolean;
  signal call_stmt_1331_call_req_0 : boolean;
  signal call_stmt_1358_call_ack_1 : boolean;
  signal call_stmt_1358_call_req_1 : boolean;
  signal RPIPE_Block1_done_1349_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1339_inst_ack_1 : boolean;
  signal RPIPE_Block1_done_1349_inst_req_0 : boolean;
  signal WPIPE_Block2_start_1339_inst_req_1 : boolean;
  signal call_stmt_1358_call_ack_0 : boolean;
  signal call_stmt_1358_call_req_0 : boolean;
  signal RPIPE_Block3_done_1355_inst_ack_1 : boolean;
  signal WPIPE_Block2_start_1339_inst_ack_0 : boolean;
  signal WPIPE_Block2_start_1339_inst_req_0 : boolean;
  signal WPIPE_Block1_start_1336_inst_req_1 : boolean;
  signal WPIPE_Block0_start_1333_inst_req_1 : boolean;
  signal RPIPE_Block0_done_1346_inst_ack_1 : boolean;
  signal WPIPE_Block1_start_1336_inst_ack_0 : boolean;
  signal RPIPE_Block2_done_1352_inst_ack_1 : boolean;
  signal RPIPE_Block3_done_1355_inst_req_1 : boolean;
  signal RPIPE_Block2_done_1352_inst_req_1 : boolean;
  signal WPIPE_Block1_start_1336_inst_req_0 : boolean;
  signal RPIPE_Block0_done_1346_inst_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTranspose_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTranspose_CP_3910_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTranspose_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3910_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTranspose_CP_3910_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTranspose_CP_3910_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTranspose_CP_3910: Block -- control-path 
    signal convTranspose_CP_3910_elements: BooleanArray(21 downto 0);
    -- 
  begin -- 
    convTranspose_CP_3910_elements(0) <= convTranspose_CP_3910_start;
    convTranspose_CP_3910_symbol <= convTranspose_CP_3910_elements(21);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_1329/branch_block_stmt_1329__entry__
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/$entry
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1329/$entry
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331__entry__
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Update/ccr
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Sample/crr
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_update_start_
      -- CP-element group 0: 	 $entry
      -- 
    ccr_3941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(0), ack => call_stmt_1331_call_req_1); -- 
    crr_3936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(0), ack => call_stmt_1331_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_sample_completed_
      -- 
    cra_3937_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1331_call_ack_0, ack => convTranspose_CP_3910_elements(1)); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	9 
    -- CP-element group 2:  members (31) 
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1329/call_stmt_1331__exit__
      -- CP-element group 2: 	 branch_block_stmt_1329/call_stmt_1331/$exit
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356__entry__
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1329/call_stmt_1331/call_stmt_1331_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Sample/req
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Sample/req
      -- 
    cca_3942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1331_call_ack_1, ack => convTranspose_CP_3910_elements(2)); -- 
    rr_4009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block0_done_1346_inst_req_0); -- 
    rr_4051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block3_done_1355_inst_req_0); -- 
    rr_4037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block2_done_1352_inst_req_0); -- 
    req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block0_start_1333_inst_req_0); -- 
    req_3995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block3_start_1342_inst_req_0); -- 
    rr_4023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => RPIPE_Block1_done_1349_inst_req_0); -- 
    req_3981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block2_start_1339_inst_req_0); -- 
    req_3967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(2), ack => WPIPE_Block1_start_1336_inst_req_0); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Sample/ack
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_update_start_
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Update/req
      -- 
    ack_3954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1333_inst_ack_0, ack => convTranspose_CP_3910_elements(3)); -- 
    req_3958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(3), ack => WPIPE_Block0_start_1333_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Update/ack
      -- CP-element group 4: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block0_start_1333_Update/$exit
      -- 
    ack_3959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_start_1333_inst_ack_1, ack => convTranspose_CP_3910_elements(4)); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_update_start_
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Update/req
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Sample/$exit
      -- 
    ack_3968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1336_inst_ack_0, ack => convTranspose_CP_3910_elements(5)); -- 
    req_3972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(5), ack => WPIPE_Block1_start_1336_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	19 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Update/ack
      -- CP-element group 6: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block1_start_1336_Update/$exit
      -- 
    ack_3973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_start_1336_inst_ack_1, ack => convTranspose_CP_3910_elements(6)); -- 
    -- CP-element group 7:  transition  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (6) 
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Update/req
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Sample/ack
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_update_start_
      -- 
    ack_3982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1339_inst_ack_0, ack => convTranspose_CP_3910_elements(7)); -- 
    req_3986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(7), ack => WPIPE_Block2_start_1339_inst_req_1); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	19 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Update/ack
      -- CP-element group 8: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block2_start_1339_update_completed_
      -- 
    ack_3987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_start_1339_inst_ack_1, ack => convTranspose_CP_3910_elements(8)); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Update/req
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Sample/ack
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_update_start_
      -- CP-element group 9: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_sample_completed_
      -- 
    ack_3996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1342_inst_ack_0, ack => convTranspose_CP_3910_elements(9)); -- 
    req_4000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(9), ack => WPIPE_Block3_start_1342_inst_req_1); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	19 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Update/ack
      -- CP-element group 10: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/WPIPE_Block3_start_1342_update_completed_
      -- 
    ack_4001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_start_1342_inst_ack_1, ack => convTranspose_CP_3910_elements(10)); -- 
    -- CP-element group 11:  transition  input  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (6) 
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_update_start_
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Sample/ra
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Update/cr
      -- CP-element group 11: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Update/$entry
      -- 
    ra_4010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1346_inst_ack_0, ack => convTranspose_CP_3910_elements(11)); -- 
    cr_4014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(11), ack => RPIPE_Block0_done_1346_inst_req_1); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	19 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Update/ca
      -- CP-element group 12: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block0_done_1346_Update/$exit
      -- 
    ca_4015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_done_1346_inst_ack_1, ack => convTranspose_CP_3910_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (6) 
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Update/cr
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Sample/ra
      -- CP-element group 13: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Sample/$exit
      -- 
    ra_4024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1349_inst_ack_0, ack => convTranspose_CP_3910_elements(13)); -- 
    cr_4028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(13), ack => RPIPE_Block1_done_1349_inst_req_1); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	19 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block1_done_1349_Update/$exit
      -- 
    ca_4029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_done_1349_inst_ack_1, ack => convTranspose_CP_3910_elements(14)); -- 
    -- CP-element group 15:  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_update_start_
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Update/cr
      -- CP-element group 15: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Update/$entry
      -- 
    ra_4038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1352_inst_ack_0, ack => convTranspose_CP_3910_elements(15)); -- 
    cr_4042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(15), ack => RPIPE_Block2_done_1352_inst_req_1); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	19 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block2_done_1352_Update/$exit
      -- 
    ca_4043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_done_1352_inst_ack_1, ack => convTranspose_CP_3910_elements(16)); -- 
    -- CP-element group 17:  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Update/cr
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Update/$entry
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_update_start_
      -- CP-element group 17: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_sample_completed_
      -- 
    ra_4052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1355_inst_ack_0, ack => convTranspose_CP_3910_elements(17)); -- 
    cr_4056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(17), ack => RPIPE_Block3_done_1355_inst_req_1); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/RPIPE_Block3_done_1355_update_completed_
      -- 
    ca_4057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_done_1355_inst_ack_1, ack => convTranspose_CP_3910_elements(18)); -- 
    -- CP-element group 19:  join  fork  transition  place  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: 	12 
    -- CP-element group 19: 	6 
    -- CP-element group 19: 	4 
    -- CP-element group 19: 	8 
    -- CP-element group 19: 	16 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	14 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19:  members (10) 
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358__entry__
      -- CP-element group 19: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356__exit__
      -- CP-element group 19: 	 branch_block_stmt_1329/assign_stmt_1335_to_assign_stmt_1356/$exit
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Update/ccr
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Update/$entry
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Sample/crr
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Sample/$entry
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_update_start_
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_sample_start_
      -- CP-element group 19: 	 branch_block_stmt_1329/call_stmt_1358/$entry
      -- 
    ccr_4073_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_4073_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(19), ack => call_stmt_1358_call_req_1); -- 
    crr_4068_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_4068_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTranspose_CP_3910_elements(19), ack => call_stmt_1358_call_req_0); -- 
    convTranspose_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 33) := "convTranspose_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= convTranspose_CP_3910_elements(10) & convTranspose_CP_3910_elements(12) & convTranspose_CP_3910_elements(6) & convTranspose_CP_3910_elements(4) & convTranspose_CP_3910_elements(8) & convTranspose_CP_3910_elements(16) & convTranspose_CP_3910_elements(18) & convTranspose_CP_3910_elements(14);
      gj_convTranspose_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTranspose_CP_3910_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Sample/cra
      -- CP-element group 20: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_sample_completed_
      -- 
    cra_4069_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_0, ack => convTranspose_CP_3910_elements(20)); -- 
    -- CP-element group 21:  transition  place  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (16) 
      -- CP-element group 21: 	 branch_block_stmt_1329/merge_stmt_1360_PhiAck/$entry
      -- CP-element group 21: 	 branch_block_stmt_1329/merge_stmt_1360_PhiAck/$exit
      -- CP-element group 21: 	 branch_block_stmt_1329/merge_stmt_1360__exit__
      -- CP-element group 21: 	 branch_block_stmt_1329/$exit
      -- CP-element group 21: 	 branch_block_stmt_1329/return__
      -- CP-element group 21: 	 branch_block_stmt_1329/return___PhiReq/$exit
      -- CP-element group 21: 	 branch_block_stmt_1329/call_stmt_1358__exit__
      -- CP-element group 21: 	 branch_block_stmt_1329/branch_block_stmt_1329__exit__
      -- CP-element group 21: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Update/cca
      -- CP-element group 21: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_1329/merge_stmt_1360_PhiReqMerge
      -- CP-element group 21: 	 branch_block_stmt_1329/call_stmt_1358/call_stmt_1358_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1329/call_stmt_1358/$exit
      -- CP-element group 21: 	 branch_block_stmt_1329/return___PhiReq/$entry
      -- CP-element group 21: 	 $exit
      -- CP-element group 21: 	 branch_block_stmt_1329/merge_stmt_1360_PhiAck/dummy
      -- 
    cca_4074_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_1, ack => convTranspose_CP_3910_elements(21)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal call11_1356 : std_logic_vector(15 downto 0);
    signal call5_1347 : std_logic_vector(15 downto 0);
    signal call7_1350 : std_logic_vector(15 downto 0);
    signal call9_1353 : std_logic_vector(15 downto 0);
    signal call_1331 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    -- shared inport operator group (0) : RPIPE_Block0_done_1346_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_done_1346_inst_req_0;
      RPIPE_Block0_done_1346_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_done_1346_inst_req_1;
      RPIPE_Block0_done_1346_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call5_1347 <= data_out(15 downto 0);
      Block0_done_read_0_gI: SplitGuardInterface generic map(name => "Block0_done_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_done_read_0: InputPortRevised -- 
        generic map ( name => "Block0_done_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_done_pipe_read_req(0),
          oack => Block0_done_pipe_read_ack(0),
          odata => Block0_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_Block1_done_1349_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_done_1349_inst_req_0;
      RPIPE_Block1_done_1349_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_done_1349_inst_req_1;
      RPIPE_Block1_done_1349_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call7_1350 <= data_out(15 downto 0);
      Block1_done_read_1_gI: SplitGuardInterface generic map(name => "Block1_done_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_done_read_1: InputPortRevised -- 
        generic map ( name => "Block1_done_read_1", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_done_pipe_read_req(0),
          oack => Block1_done_pipe_read_ack(0),
          odata => Block1_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_Block2_done_1352_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_done_1352_inst_req_0;
      RPIPE_Block2_done_1352_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_done_1352_inst_req_1;
      RPIPE_Block2_done_1352_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call9_1353 <= data_out(15 downto 0);
      Block2_done_read_2_gI: SplitGuardInterface generic map(name => "Block2_done_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_done_read_2: InputPortRevised -- 
        generic map ( name => "Block2_done_read_2", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_done_pipe_read_req(0),
          oack => Block2_done_pipe_read_ack(0),
          odata => Block2_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : RPIPE_Block3_done_1355_inst 
    InportGroup_3: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_done_1355_inst_req_0;
      RPIPE_Block3_done_1355_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_done_1355_inst_req_1;
      RPIPE_Block3_done_1355_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call11_1356 <= data_out(15 downto 0);
      Block3_done_read_3_gI: SplitGuardInterface generic map(name => "Block3_done_read_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_done_read_3: InputPortRevised -- 
        generic map ( name => "Block3_done_read_3", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_done_pipe_read_req(0),
          oack => Block3_done_pipe_read_ack(0),
          odata => Block3_done_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : WPIPE_Block0_start_1333_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_start_1333_inst_req_0;
      WPIPE_Block0_start_1333_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_start_1333_inst_req_1;
      WPIPE_Block0_start_1333_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1331;
      Block0_start_write_0_gI: SplitGuardInterface generic map(name => "Block0_start_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_start_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_start_pipe_write_req(0),
          oack => Block0_start_pipe_write_ack(0),
          odata => Block0_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_Block1_start_1336_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_start_1336_inst_req_0;
      WPIPE_Block1_start_1336_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_start_1336_inst_req_1;
      WPIPE_Block1_start_1336_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1331;
      Block1_start_write_1_gI: SplitGuardInterface generic map(name => "Block1_start_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_start_write_1: OutputPortRevised -- 
        generic map ( name => "Block1_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_start_pipe_write_req(0),
          oack => Block1_start_pipe_write_ack(0),
          odata => Block1_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_Block2_start_1339_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_start_1339_inst_req_0;
      WPIPE_Block2_start_1339_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_start_1339_inst_req_1;
      WPIPE_Block2_start_1339_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1331;
      Block2_start_write_2_gI: SplitGuardInterface generic map(name => "Block2_start_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_start_write_2: OutputPortRevised -- 
        generic map ( name => "Block2_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_start_pipe_write_req(0),
          oack => Block2_start_pipe_write_ack(0),
          odata => Block2_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_Block3_start_1342_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_start_1342_inst_req_0;
      WPIPE_Block3_start_1342_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_start_1342_inst_req_1;
      WPIPE_Block3_start_1342_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1331;
      Block3_start_write_3_gI: SplitGuardInterface generic map(name => "Block3_start_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_start_write_3: OutputPortRevised -- 
        generic map ( name => "Block3_start", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_start_pipe_write_req(0),
          oack => Block3_start_pipe_write_ack(0),
          odata => Block3_start_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared call operator group (0) : call_stmt_1331_call 
    testConfigure_call_group_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1331_call_req_0;
      call_stmt_1331_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1331_call_req_1;
      call_stmt_1331_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      testConfigure_call_group_0_gI: SplitGuardInterface generic map(name => "testConfigure_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      call_1331 <= data_out(15 downto 0);
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => testConfigure_call_reqs(0),
          ackR => testConfigure_call_acks(0),
          tagR => testConfigure_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 16,
          owidth => 16,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => testConfigure_return_acks(0), -- cross-over
          ackL => testConfigure_return_reqs(0), -- cross-over
          dataL => testConfigure_return_data(15 downto 0),
          tagL => testConfigure_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1358_call 
    sendOutput_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1358_call_req_0;
      call_stmt_1358_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1358_call_req_1;
      call_stmt_1358_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      sendOutput_call_group_1_gI: SplitGuardInterface generic map(name => "sendOutput_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (name => "InputMuxBaseNoData",
        twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendOutput_call_reqs(0),
          ackR => sendOutput_call_acks(0),
          tagR => sendOutput_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendOutput_return_acks(0), -- cross-over
          ackL => sendOutput_return_reqs(0), -- cross-over
          tagL => sendOutput_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end convTranspose_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeA is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeA;
architecture convTransposeA_arch of convTransposeA is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeA_CP_4083_start: Boolean;
  signal convTransposeA_CP_4083_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1690_load_0_req_1 : boolean;
  signal addr_of_1686_final_reg_req_0 : boolean;
  signal type_cast_1679_inst_req_1 : boolean;
  signal ptr_deref_1690_load_0_ack_1 : boolean;
  signal ptr_deref_1492_load_0_ack_0 : boolean;
  signal type_cast_1679_inst_ack_1 : boolean;
  signal addr_of_1686_final_reg_ack_0 : boolean;
  signal array_obj_ref_1716_index_offset_req_0 : boolean;
  signal ptr_deref_1690_load_0_ack_0 : boolean;
  signal ptr_deref_1492_load_0_req_0 : boolean;
  signal addr_of_1717_final_reg_req_0 : boolean;
  signal addr_of_1717_final_reg_ack_0 : boolean;
  signal type_cast_1710_inst_ack_1 : boolean;
  signal type_cast_1710_inst_req_1 : boolean;
  signal array_obj_ref_1716_index_offset_ack_1 : boolean;
  signal array_obj_ref_1716_index_offset_req_1 : boolean;
  signal type_cast_1710_inst_req_0 : boolean;
  signal type_cast_1710_inst_ack_0 : boolean;
  signal type_cast_1521_inst_req_0 : boolean;
  signal ptr_deref_1690_load_0_req_0 : boolean;
  signal type_cast_1679_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1366_inst_req_0 : boolean;
  signal RPIPE_Block0_start_1366_inst_ack_0 : boolean;
  signal RPIPE_Block0_start_1366_inst_req_1 : boolean;
  signal RPIPE_Block0_start_1366_inst_ack_1 : boolean;
  signal array_obj_ref_1685_index_offset_ack_1 : boolean;
  signal type_cast_1679_inst_req_0 : boolean;
  signal array_obj_ref_1685_index_offset_req_1 : boolean;
  signal type_cast_1648_inst_ack_1 : boolean;
  signal ptr_deref_1474_load_0_ack_1 : boolean;
  signal type_cast_1648_inst_req_1 : boolean;
  signal array_obj_ref_1685_index_offset_ack_0 : boolean;
  signal ptr_deref_1379_load_0_req_0 : boolean;
  signal ptr_deref_1379_load_0_ack_0 : boolean;
  signal ptr_deref_1474_load_0_req_1 : boolean;
  signal array_obj_ref_1685_index_offset_req_0 : boolean;
  signal ptr_deref_1379_load_0_req_1 : boolean;
  signal ptr_deref_1379_load_0_ack_1 : boolean;
  signal type_cast_1648_inst_ack_0 : boolean;
  signal type_cast_1648_inst_req_0 : boolean;
  signal ptr_deref_1391_load_0_req_0 : boolean;
  signal type_cast_1526_inst_ack_1 : boolean;
  signal ptr_deref_1391_load_0_ack_0 : boolean;
  signal ptr_deref_1391_load_0_req_1 : boolean;
  signal type_cast_1526_inst_req_1 : boolean;
  signal ptr_deref_1391_load_0_ack_1 : boolean;
  signal addr_of_1686_final_reg_ack_1 : boolean;
  signal type_cast_1526_inst_ack_0 : boolean;
  signal type_cast_1526_inst_req_0 : boolean;
  signal type_cast_1521_inst_ack_1 : boolean;
  signal type_cast_1521_inst_req_1 : boolean;
  signal ptr_deref_1492_load_0_ack_1 : boolean;
  signal ptr_deref_1401_load_0_req_0 : boolean;
  signal ptr_deref_1401_load_0_ack_0 : boolean;
  signal ptr_deref_1492_load_0_req_1 : boolean;
  signal ptr_deref_1401_load_0_req_1 : boolean;
  signal ptr_deref_1401_load_0_ack_1 : boolean;
  signal type_cast_1521_inst_ack_0 : boolean;
  signal addr_of_1686_final_reg_req_1 : boolean;
  signal type_cast_1405_inst_req_0 : boolean;
  signal type_cast_1405_inst_ack_0 : boolean;
  signal type_cast_1405_inst_req_1 : boolean;
  signal type_cast_1405_inst_ack_1 : boolean;
  signal ptr_deref_1417_load_0_req_0 : boolean;
  signal ptr_deref_1417_load_0_ack_0 : boolean;
  signal ptr_deref_1417_load_0_req_1 : boolean;
  signal ptr_deref_1417_load_0_ack_1 : boolean;
  signal LOAD_padding_1420_load_0_req_0 : boolean;
  signal LOAD_padding_1420_load_0_ack_0 : boolean;
  signal array_obj_ref_1716_index_offset_ack_0 : boolean;
  signal LOAD_padding_1420_load_0_req_1 : boolean;
  signal LOAD_padding_1420_load_0_ack_1 : boolean;
  signal type_cast_1424_inst_req_0 : boolean;
  signal type_cast_1424_inst_ack_0 : boolean;
  signal type_cast_1424_inst_req_1 : boolean;
  signal type_cast_1424_inst_ack_1 : boolean;
  signal ptr_deref_1434_load_0_req_0 : boolean;
  signal ptr_deref_1434_load_0_ack_0 : boolean;
  signal ptr_deref_1434_load_0_req_1 : boolean;
  signal ptr_deref_1434_load_0_ack_1 : boolean;
  signal type_cast_1438_inst_req_0 : boolean;
  signal type_cast_1438_inst_ack_0 : boolean;
  signal type_cast_1438_inst_req_1 : boolean;
  signal type_cast_1438_inst_ack_1 : boolean;
  signal ptr_deref_1450_load_0_req_0 : boolean;
  signal ptr_deref_1450_load_0_ack_0 : boolean;
  signal ptr_deref_1450_load_0_req_1 : boolean;
  signal ptr_deref_1450_load_0_ack_1 : boolean;
  signal ptr_deref_1462_load_0_req_0 : boolean;
  signal ptr_deref_1462_load_0_ack_0 : boolean;
  signal ptr_deref_1462_load_0_req_1 : boolean;
  signal ptr_deref_1462_load_0_ack_1 : boolean;
  signal ptr_deref_1474_load_0_req_0 : boolean;
  signal ptr_deref_1474_load_0_ack_0 : boolean;
  signal addr_of_1717_final_reg_req_1 : boolean;
  signal addr_of_1717_final_reg_ack_1 : boolean;
  signal ptr_deref_1720_store_0_req_0 : boolean;
  signal ptr_deref_1720_store_0_ack_0 : boolean;
  signal ptr_deref_1720_store_0_req_1 : boolean;
  signal ptr_deref_1720_store_0_ack_1 : boolean;
  signal type_cast_1726_inst_req_0 : boolean;
  signal type_cast_1726_inst_ack_0 : boolean;
  signal type_cast_1726_inst_req_1 : boolean;
  signal type_cast_1726_inst_ack_1 : boolean;
  signal if_stmt_1739_branch_req_0 : boolean;
  signal if_stmt_1739_branch_ack_1 : boolean;
  signal if_stmt_1739_branch_ack_0 : boolean;
  signal type_cast_1763_inst_req_0 : boolean;
  signal type_cast_1763_inst_ack_0 : boolean;
  signal type_cast_1763_inst_req_1 : boolean;
  signal type_cast_1763_inst_ack_1 : boolean;
  signal type_cast_1772_inst_req_0 : boolean;
  signal type_cast_1772_inst_ack_0 : boolean;
  signal type_cast_1772_inst_req_1 : boolean;
  signal type_cast_1772_inst_ack_1 : boolean;
  signal type_cast_1789_inst_req_0 : boolean;
  signal type_cast_1789_inst_ack_0 : boolean;
  signal type_cast_1789_inst_req_1 : boolean;
  signal type_cast_1789_inst_ack_1 : boolean;
  signal if_stmt_1796_branch_req_0 : boolean;
  signal if_stmt_1796_branch_ack_1 : boolean;
  signal if_stmt_1796_branch_ack_0 : boolean;
  signal WPIPE_Block0_done_1804_inst_req_0 : boolean;
  signal WPIPE_Block0_done_1804_inst_ack_0 : boolean;
  signal WPIPE_Block0_done_1804_inst_req_1 : boolean;
  signal WPIPE_Block0_done_1804_inst_ack_1 : boolean;
  signal phi_stmt_1502_req_0 : boolean;
  signal phi_stmt_1509_req_0 : boolean;
  signal type_cast_1508_inst_req_0 : boolean;
  signal type_cast_1508_inst_ack_0 : boolean;
  signal type_cast_1508_inst_req_1 : boolean;
  signal type_cast_1508_inst_ack_1 : boolean;
  signal phi_stmt_1502_req_1 : boolean;
  signal type_cast_1515_inst_req_0 : boolean;
  signal type_cast_1515_inst_ack_0 : boolean;
  signal type_cast_1515_inst_req_1 : boolean;
  signal type_cast_1515_inst_ack_1 : boolean;
  signal phi_stmt_1509_req_1 : boolean;
  signal phi_stmt_1502_ack_0 : boolean;
  signal phi_stmt_1509_ack_0 : boolean;
  signal type_cast_1638_inst_req_0 : boolean;
  signal type_cast_1638_inst_ack_0 : boolean;
  signal type_cast_1638_inst_req_1 : boolean;
  signal type_cast_1638_inst_ack_1 : boolean;
  signal phi_stmt_1632_req_1 : boolean;
  signal phi_stmt_1632_req_0 : boolean;
  signal phi_stmt_1632_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeA_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeA_CP_4083_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeA_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeA_CP_4083_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeA_CP_4083: Block -- control-path 
    signal convTransposeA_CP_4083_elements: BooleanArray(88 downto 0);
    -- 
  begin -- 
    convTransposeA_CP_4083_elements(0) <= convTransposeA_CP_4083_start;
    convTransposeA_CP_4083_symbol <= convTransposeA_CP_4083_elements(68);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1364/$entry
      -- CP-element group 0: 	 branch_block_stmt_1364/branch_block_stmt_1364__entry__
      -- CP-element group 0: 	 branch_block_stmt_1364/assign_stmt_1367__entry__
      -- CP-element group 0: 	 branch_block_stmt_1364/assign_stmt_1367/$entry
      -- CP-element group 0: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Sample/rr
      -- 
    rr_4131_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4131_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(0), ack => RPIPE_Block0_start_1366_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Update/cr
      -- 
    ra_4132_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1366_inst_ack_0, ack => convTransposeA_CP_4083_elements(1)); -- 
    cr_4136_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4136_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(1), ack => RPIPE_Block0_start_1366_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	5 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2:  members (262) 
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1367__exit__
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499__entry__
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1367/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1367/RPIPE_Block0_start_1366_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/word_0/rr
      -- 
    ca_4137_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block0_start_1366_inst_ack_1, ack => convTransposeA_CP_4083_elements(2)); -- 
    rr_4648_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4648_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1492_load_0_req_0); -- 
    rr_4173_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4173_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1379_load_0_req_0); -- 
    cr_4609_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4609_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1474_load_0_req_1); -- 
    cr_4184_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4184_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1379_load_0_req_1); -- 
    rr_4223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1391_load_0_req_0); -- 
    cr_4234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1391_load_0_req_1); -- 
    rr_4273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1401_load_0_req_0); -- 
    cr_4659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1492_load_0_req_1); -- 
    cr_4284_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4284_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1401_load_0_req_1); -- 
    cr_4303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1405_inst_req_1); -- 
    rr_4337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1417_load_0_req_0); -- 
    cr_4348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1417_load_0_req_1); -- 
    rr_4370_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4370_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => LOAD_padding_1420_load_0_req_0); -- 
    cr_4381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => LOAD_padding_1420_load_0_req_1); -- 
    cr_4400_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4400_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1424_inst_req_1); -- 
    rr_4434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1434_load_0_req_0); -- 
    cr_4445_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4445_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1434_load_0_req_1); -- 
    cr_4464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => type_cast_1438_inst_req_1); -- 
    rr_4498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1450_load_0_req_0); -- 
    cr_4509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1450_load_0_req_1); -- 
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1462_load_0_req_0); -- 
    cr_4559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1462_load_0_req_1); -- 
    rr_4598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(2), ack => ptr_deref_1474_load_0_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Sample/word_access_start/word_0/ra
      -- 
    ra_4174_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1379_load_0_ack_0, ack => convTransposeA_CP_4083_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	29 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/ptr_deref_1379_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/ptr_deref_1379_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/ptr_deref_1379_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1379_Update/ptr_deref_1379_Merge/merge_ack
      -- 
    ca_4185_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1379_load_0_ack_1, ack => convTransposeA_CP_4083_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Sample/word_access_start/word_0/ra
      -- 
    ra_4224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1391_load_0_ack_0, ack => convTransposeA_CP_4083_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	29 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/ptr_deref_1391_Merge/$entry
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/ptr_deref_1391_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/ptr_deref_1391_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1391_Update/ptr_deref_1391_Merge/merge_ack
      -- 
    ca_4235_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1391_load_0_ack_1, ack => convTransposeA_CP_4083_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Sample/word_access_start/word_0/ra
      -- 
    ra_4274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1401_load_0_ack_0, ack => convTransposeA_CP_4083_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/ptr_deref_1401_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/ptr_deref_1401_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/ptr_deref_1401_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1401_Update/ptr_deref_1401_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Sample/rr
      -- 
    ca_4285_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1401_load_0_ack_1, ack => convTransposeA_CP_4083_elements(8)); -- 
    rr_4298_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4298_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(8), ack => type_cast_1405_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Sample/ra
      -- 
    ra_4299_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_0, ack => convTransposeA_CP_4083_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	29 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1405_Update/ca
      -- 
    ca_4304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1405_inst_ack_1, ack => convTransposeA_CP_4083_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Sample/word_access_start/word_0/ra
      -- 
    ra_4338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1417_load_0_ack_0, ack => convTransposeA_CP_4083_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/ptr_deref_1417_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/ptr_deref_1417_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/ptr_deref_1417_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1417_Update/ptr_deref_1417_Merge/merge_ack
      -- 
    ca_4349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1417_load_0_ack_1, ack => convTransposeA_CP_4083_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Sample/word_access_start/word_0/ra
      -- 
    ra_4371_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1420_load_0_ack_0, ack => convTransposeA_CP_4083_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/LOAD_padding_1420_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/LOAD_padding_1420_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/LOAD_padding_1420_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/LOAD_padding_1420_Update/LOAD_padding_1420_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Sample/rr
      -- 
    ca_4382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1420_load_0_ack_1, ack => convTransposeA_CP_4083_elements(14)); -- 
    rr_4395_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4395_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(14), ack => type_cast_1424_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Sample/ra
      -- 
    ra_4396_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1424_inst_ack_0, ack => convTransposeA_CP_4083_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	29 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1424_Update/ca
      -- 
    ca_4401_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1424_inst_ack_1, ack => convTransposeA_CP_4083_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Sample/word_access_start/word_0/ra
      -- 
    ra_4435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1434_load_0_ack_0, ack => convTransposeA_CP_4083_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/ptr_deref_1434_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/ptr_deref_1434_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/ptr_deref_1434_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1434_Update/ptr_deref_1434_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Sample/rr
      -- 
    ca_4446_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1434_load_0_ack_1, ack => convTransposeA_CP_4083_elements(18)); -- 
    rr_4459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(18), ack => type_cast_1438_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Sample/ra
      -- 
    ra_4460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_0, ack => convTransposeA_CP_4083_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	29 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/type_cast_1438_Update/ca
      -- 
    ca_4465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_1, ack => convTransposeA_CP_4083_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Sample/word_access_start/word_0/ra
      -- 
    ra_4499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1450_load_0_ack_0, ack => convTransposeA_CP_4083_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	29 
    -- CP-element group 22:  members (9) 
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/ptr_deref_1450_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/ptr_deref_1450_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/ptr_deref_1450_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1450_Update/ptr_deref_1450_Merge/merge_ack
      -- 
    ca_4510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1450_load_0_ack_1, ack => convTransposeA_CP_4083_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Sample/word_access_start/word_0/ra
      -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1462_load_0_ack_0, ack => convTransposeA_CP_4083_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	29 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/ptr_deref_1462_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/ptr_deref_1462_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/ptr_deref_1462_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1462_Update/ptr_deref_1462_Merge/merge_ack
      -- 
    ca_4560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1462_load_0_ack_1, ack => convTransposeA_CP_4083_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Sample/word_access_start/word_0/ra
      -- 
    ra_4599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1474_load_0_ack_0, ack => convTransposeA_CP_4083_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	29 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/ptr_deref_1474_Merge/merge_ack
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/ptr_deref_1474_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/ptr_deref_1474_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/ptr_deref_1474_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1474_update_completed_
      -- 
    ca_4610_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1474_load_0_ack_1, ack => convTransposeA_CP_4083_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/word_0/ra
      -- CP-element group 27: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Sample/$exit
      -- 
    ra_4649_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1492_load_0_ack_0, ack => convTransposeA_CP_4083_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/ptr_deref_1492_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/ptr_deref_1492_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/ptr_deref_1492_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/ptr_deref_1492_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/ptr_deref_1492_Update/word_access_complete/word_0/ca
      -- 
    ca_4660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1492_load_0_ack_1, ack => convTransposeA_CP_4083_elements(28)); -- 
    -- CP-element group 29:  join  fork  transition  place  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	16 
    -- CP-element group 29: 	22 
    -- CP-element group 29: 	24 
    -- CP-element group 29: 	26 
    -- CP-element group 29: 	28 
    -- CP-element group 29: 	20 
    -- CP-element group 29: 	4 
    -- CP-element group 29: 	6 
    -- CP-element group 29: 	10 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	69 
    -- CP-element group 29: 	70 
    -- CP-element group 29:  members (8) 
      -- CP-element group 29: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499__exit__
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter
      -- CP-element group 29: 	 branch_block_stmt_1364/assign_stmt_1376_to_assign_stmt_1499/$exit
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/$entry
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/$entry
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/$entry
      -- CP-element group 29: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/$entry
      -- 
    convTransposeA_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(16) & convTransposeA_CP_4083_elements(22) & convTransposeA_CP_4083_elements(24) & convTransposeA_CP_4083_elements(26) & convTransposeA_CP_4083_elements(28) & convTransposeA_CP_4083_elements(20) & convTransposeA_CP_4083_elements(4) & convTransposeA_CP_4083_elements(6) & convTransposeA_CP_4083_elements(10) & convTransposeA_CP_4083_elements(12);
      gj_convTransposeA_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	82 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Sample/ra
      -- 
    ra_4677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_0, ack => convTransposeA_CP_4083_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	82 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	34 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Update/$exit
      -- 
    ca_4682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1521_inst_ack_1, ack => convTransposeA_CP_4083_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	82 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Sample/ra
      -- CP-element group 32: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_sample_completed_
      -- 
    ra_4691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_0, ack => convTransposeA_CP_4083_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	82 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_update_completed_
      -- 
    ca_4696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1526_inst_ack_1, ack => convTransposeA_CP_4083_elements(33)); -- 
    -- CP-element group 34:  join  transition  place  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	31 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	86 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629__exit__
      -- CP-element group 34: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 34: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/$exit
      -- CP-element group 34: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 34: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/$entry
      -- CP-element group 34: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$entry
      -- 
    convTransposeA_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(31) & convTransposeA_CP_4083_elements(33);
      gj_convTransposeA_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Sample/ra
      -- CP-element group 35: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_sample_completed_
      -- 
    ra_4708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_0, ack => convTransposeA_CP_4083_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	88 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	45 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (9) 
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Sample/rr
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Update/ca
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_sample_start_
      -- 
    ca_4713_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1648_inst_ack_1, ack => convTransposeA_CP_4083_elements(36)); -- 
    rr_4831_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4831_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(36), ack => type_cast_1710_inst_req_0); -- 
    rr_4721_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4721_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(36), ack => type_cast_1679_inst_req_0); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Sample/ra
      -- CP-element group 37: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_sample_completed_
      -- 
    ra_4722_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1679_inst_ack_0, ack => convTransposeA_CP_4083_elements(37)); -- 
    -- CP-element group 38:  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	88 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (16) 
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_resize_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_resize_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_computed_1
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_resized_1
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_scaled_1
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_resize_1/index_resize_req
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Sample/req
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_scale_1/scale_rename_ack
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_scale_1/scale_rename_req
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_scale_1/$exit
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_scale_1/$entry
      -- CP-element group 38: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_index_resize_1/index_resize_ack
      -- 
    ca_4727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1679_inst_ack_1, ack => convTransposeA_CP_4083_elements(38)); -- 
    req_4752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(38), ack => array_obj_ref_1685_index_offset_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	56 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Sample/ack
      -- CP-element group 39: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_sample_complete
      -- 
    ack_4753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1685_index_offset_ack_0, ack => convTransposeA_CP_4083_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	88 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (11) 
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_request/req
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_offset_calculated
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_base_plus_offset/sum_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_request/$entry
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_base_plus_offset/sum_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_base_plus_offset/$exit
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_base_plus_offset/$entry
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_root_address_calculated
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Update/ack
      -- CP-element group 40: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Update/$exit
      -- 
    ack_4758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1685_index_offset_ack_1, ack => convTransposeA_CP_4083_elements(40)); -- 
    req_4767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(40), ack => addr_of_1686_final_reg_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_request/ack
      -- CP-element group 41: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_request/$exit
      -- 
    ack_4768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1686_final_reg_ack_0, ack => convTransposeA_CP_4083_elements(41)); -- 
    -- CP-element group 42:  join  fork  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	88 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (24) 
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_complete/$exit
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_word_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_addr_resize/$entry
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_addr_resize/$exit
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_addr_resize/base_resize_req
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_word_addrgen/$entry
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_word_addrgen/root_register_ack
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_addr_resize/base_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_address_resized
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/word_0/rr
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/word_0/$entry
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_word_addrgen/root_register_req
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_complete/ack
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_word_addrgen/$exit
      -- CP-element group 42: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/$entry
      -- 
    ack_4773_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1686_final_reg_ack_1, ack => convTransposeA_CP_4083_elements(42)); -- 
    rr_4806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(42), ack => ptr_deref_1690_load_0_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (5) 
      -- CP-element group 43: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/word_0/ra
      -- CP-element group 43: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/word_0/$exit
      -- CP-element group 43: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Sample/word_access_start/$exit
      -- 
    ra_4807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1690_load_0_ack_0, ack => convTransposeA_CP_4083_elements(43)); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	88 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	51 
    -- CP-element group 44:  members (9) 
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/word_0/$exit
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/word_0/ca
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/ptr_deref_1690_Merge/merge_req
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/ptr_deref_1690_Merge/$entry
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/ptr_deref_1690_Merge/$exit
      -- CP-element group 44: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/ptr_deref_1690_Merge/merge_ack
      -- 
    ca_4818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1690_load_0_ack_1, ack => convTransposeA_CP_4083_elements(44)); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	36 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Sample/ra
      -- CP-element group 45: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_sample_completed_
      -- 
    ra_4832_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_0, ack => convTransposeA_CP_4083_elements(45)); -- 
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	88 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (16) 
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_scale_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_scale_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_resized_1
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Sample/req
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_scaled_1
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Update/ca
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_computed_1
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_scale_1/scale_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_resize_1/$entry
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_resize_1/$exit
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_resize_1/index_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_scale_1/scale_rename_req
      -- CP-element group 46: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_index_resize_1/index_resize_req
      -- 
    ca_4837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1710_inst_ack_1, ack => convTransposeA_CP_4083_elements(46)); -- 
    req_4862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(46), ack => array_obj_ref_1716_index_offset_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	56 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_sample_complete
      -- CP-element group 47: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Sample/ack
      -- 
    ack_4863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1716_index_offset_ack_0, ack => convTransposeA_CP_4083_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	88 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (11) 
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_base_plus_offset/$exit
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_base_plus_offset/sum_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_request/req
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_base_plus_offset/sum_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_base_plus_offset/$entry
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_root_address_calculated
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_offset_calculated
      -- CP-element group 48: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_request/$entry
      -- 
    ack_4868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1716_index_offset_ack_1, ack => convTransposeA_CP_4083_elements(48)); -- 
    req_4877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(48), ack => addr_of_1717_final_reg_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_request/$exit
      -- CP-element group 49: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_request/ack
      -- CP-element group 49: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_sample_completed_
      -- 
    ack_4878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1717_final_reg_ack_0, ack => convTransposeA_CP_4083_elements(49)); -- 
    -- CP-element group 50:  fork  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	88 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (19) 
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_complete/ack
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_word_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_address_resized
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_addr_resize/$entry
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_addr_resize/$exit
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_addr_resize/base_resize_req
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_addr_resize/base_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_word_addrgen/$entry
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_word_addrgen/$exit
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_word_addrgen/root_register_req
      -- CP-element group 50: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_word_addrgen/root_register_ack
      -- 
    ack_4883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1717_final_reg_ack_1, ack => convTransposeA_CP_4083_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	44 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (9) 
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/ptr_deref_1720_Split/$entry
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/ptr_deref_1720_Split/$exit
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/ptr_deref_1720_Split/split_req
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/ptr_deref_1720_Split/split_ack
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/word_0/rr
      -- 
    rr_4921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(51), ack => ptr_deref_1720_store_0_req_0); -- 
    convTransposeA_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(44) & convTransposeA_CP_4083_elements(50);
      gj_convTransposeA_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Sample/word_access_start/word_0/ra
      -- 
    ra_4922_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_store_0_ack_0, ack => convTransposeA_CP_4083_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	88 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	56 
    -- CP-element group 53:  members (5) 
      -- CP-element group 53: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/word_0/ca
      -- 
    ca_4933_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1720_store_0_ack_1, ack => convTransposeA_CP_4083_elements(53)); -- 
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	88 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Sample/ra
      -- 
    ra_4942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1726_inst_ack_0, ack => convTransposeA_CP_4083_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	88 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Update/ca
      -- 
    ca_4947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1726_inst_ack_1, ack => convTransposeA_CP_4083_elements(55)); -- 
    -- CP-element group 56:  branch  join  transition  place  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	47 
    -- CP-element group 56: 	53 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	39 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (10) 
      -- CP-element group 56: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738__exit__
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739__entry__
      -- CP-element group 56: 	 branch_block_stmt_1364/R_cmp_1740_place
      -- CP-element group 56: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/$exit
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_dead_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_eval_test/$entry
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_eval_test/$exit
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_eval_test/branch_req
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_if_link/$entry
      -- CP-element group 56: 	 branch_block_stmt_1364/if_stmt_1739_else_link/$entry
      -- 
    branch_req_4955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_4955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(56), ack => if_stmt_1739_branch_req_0); -- 
    convTransposeA_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(47) & convTransposeA_CP_4083_elements(53) & convTransposeA_CP_4083_elements(55) & convTransposeA_CP_4083_elements(39);
      gj_convTransposeA_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	83 
    -- CP-element group 57: 	84 
    -- CP-element group 57:  members (24) 
      -- CP-element group 57: 	 branch_block_stmt_1364/whilex_xbody_ifx_xthen
      -- CP-element group 57: 	 branch_block_stmt_1364/merge_stmt_1745__exit__
      -- CP-element group 57: 	 branch_block_stmt_1364/assign_stmt_1751__entry__
      -- CP-element group 57: 	 branch_block_stmt_1364/assign_stmt_1751__exit__
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody
      -- CP-element group 57: 	 branch_block_stmt_1364/if_stmt_1739_if_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_1364/if_stmt_1739_if_link/if_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_1364/assign_stmt_1751/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/assign_stmt_1751/$exit
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/rr
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/cr
      -- CP-element group 57: 	 branch_block_stmt_1364/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_1364/merge_stmt_1745_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_1364/merge_stmt_1745_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_1364/merge_stmt_1745_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_1364/merge_stmt_1745_PhiAck/dummy
      -- 
    if_choice_transition_4960_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1739_branch_ack_1, ack => convTransposeA_CP_4083_elements(57)); -- 
    rr_5143_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5143_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(57), ack => type_cast_1638_inst_req_0); -- 
    cr_5148_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5148_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(57), ack => type_cast_1638_inst_req_1); -- 
    -- CP-element group 58:  fork  transition  place  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58: 	62 
    -- CP-element group 58: 	64 
    -- CP-element group 58:  members (24) 
      -- CP-element group 58: 	 branch_block_stmt_1364/whilex_xbody_ifx_xelse
      -- CP-element group 58: 	 branch_block_stmt_1364/merge_stmt_1753__exit__
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795__entry__
      -- CP-element group 58: 	 branch_block_stmt_1364/if_stmt_1739_else_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1364/if_stmt_1739_else_link/else_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Sample/rr
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_update_start_
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Update/cr
      -- CP-element group 58: 	 branch_block_stmt_1364/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1364/merge_stmt_1753_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1364/merge_stmt_1753_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1364/merge_stmt_1753_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1364/merge_stmt_1753_PhiAck/dummy
      -- 
    else_choice_transition_4964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1739_branch_ack_0, ack => convTransposeA_CP_4083_elements(58)); -- 
    rr_4980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1763_inst_req_0); -- 
    cr_4985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1763_inst_req_1); -- 
    cr_4999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1772_inst_req_1); -- 
    cr_5013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(58), ack => type_cast_1789_inst_req_1); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Sample/$exit
      -- CP-element group 59: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Sample/ra
      -- 
    ra_4981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_0, ack => convTransposeA_CP_4083_elements(59)); -- 
    -- CP-element group 60:  transition  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (6) 
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1763_Update/ca
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Sample/rr
      -- 
    ca_4986_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1763_inst_ack_1, ack => convTransposeA_CP_4083_elements(60)); -- 
    rr_4994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(60), ack => type_cast_1772_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Sample/ra
      -- 
    ra_4995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_0, ack => convTransposeA_CP_4083_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	58 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1772_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Sample/rr
      -- 
    ca_5000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1772_inst_ack_1, ack => convTransposeA_CP_4083_elements(62)); -- 
    rr_5008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(62), ack => type_cast_1789_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Sample/ra
      -- 
    ra_5009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_0, ack => convTransposeA_CP_4083_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	58 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_1364/R_cmp77_1797_place
      -- CP-element group 64: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795__exit__
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796__entry__
      -- CP-element group 64: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/$exit
      -- CP-element group 64: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_1364/assign_stmt_1759_to_assign_stmt_1795/type_cast_1789_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_1364/if_stmt_1796_else_link/$entry
      -- 
    ca_5014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1789_inst_ack_1, ack => convTransposeA_CP_4083_elements(64)); -- 
    branch_req_5022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_5022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(64), ack => if_stmt_1796_branch_req_0); -- 
    -- CP-element group 65:  merge  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (15) 
      -- CP-element group 65: 	 branch_block_stmt_1364/ifx_xelse_whilex_xend
      -- CP-element group 65: 	 branch_block_stmt_1364/merge_stmt_1802__exit__
      -- CP-element group 65: 	 branch_block_stmt_1364/assign_stmt_1806__entry__
      -- CP-element group 65: 	 branch_block_stmt_1364/if_stmt_1796_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_1364/if_stmt_1796_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_1364/assign_stmt_1806/$entry
      -- CP-element group 65: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1364/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_1364/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_1364/merge_stmt_1802_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_1364/merge_stmt_1802_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_1364/merge_stmt_1802_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1364/merge_stmt_1802_PhiAck/dummy
      -- 
    if_choice_transition_5027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1796_branch_ack_1, ack => convTransposeA_CP_4083_elements(65)); -- 
    req_5044_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5044_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(65), ack => WPIPE_Block0_done_1804_inst_req_0); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	72 
    -- CP-element group 66: 	73 
    -- CP-element group 66: 	75 
    -- CP-element group 66: 	76 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 66: 	 branch_block_stmt_1364/if_stmt_1796_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_1364/if_stmt_1796_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Update/cr
      -- 
    else_choice_transition_5031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1796_branch_ack_0, ack => convTransposeA_CP_4083_elements(66)); -- 
    rr_5088_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5088_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1508_inst_req_0); -- 
    cr_5093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1508_inst_req_1); -- 
    rr_5111_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5111_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1515_inst_req_0); -- 
    cr_5116_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5116_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(66), ack => type_cast_1515_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Sample/ack
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Update/req
      -- 
    ack_5045_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1804_inst_ack_0, ack => convTransposeA_CP_4083_elements(67)); -- 
    req_5049_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5049_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(67), ack => WPIPE_Block0_done_1804_inst_req_1); -- 
    -- CP-element group 68:  transition  place  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (16) 
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 branch_block_stmt_1364/$exit
      -- CP-element group 68: 	 branch_block_stmt_1364/branch_block_stmt_1364__exit__
      -- CP-element group 68: 	 branch_block_stmt_1364/assign_stmt_1806__exit__
      -- CP-element group 68: 	 branch_block_stmt_1364/return__
      -- CP-element group 68: 	 branch_block_stmt_1364/merge_stmt_1808__exit__
      -- CP-element group 68: 	 branch_block_stmt_1364/assign_stmt_1806/$exit
      -- CP-element group 68: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1364/assign_stmt_1806/WPIPE_Block0_done_1804_Update/ack
      -- CP-element group 68: 	 branch_block_stmt_1364/return___PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_1364/return___PhiReq/$exit
      -- CP-element group 68: 	 branch_block_stmt_1364/merge_stmt_1808_PhiReqMerge
      -- CP-element group 68: 	 branch_block_stmt_1364/merge_stmt_1808_PhiAck/$entry
      -- CP-element group 68: 	 branch_block_stmt_1364/merge_stmt_1808_PhiAck/$exit
      -- CP-element group 68: 	 branch_block_stmt_1364/merge_stmt_1808_PhiAck/dummy
      -- 
    ack_5050_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block0_done_1804_inst_ack_1, ack => convTransposeA_CP_4083_elements(68)); -- 
    -- CP-element group 69:  transition  output  delay-element  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	29 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/$exit
      -- CP-element group 69: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/$exit
      -- CP-element group 69: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1506_konst_delay_trans
      -- CP-element group 69: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_req
      -- 
    phi_stmt_1502_req_5061_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1502_req_5061_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(69), ack => phi_stmt_1502_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(69) is a control-delay.
    cp_element_69_delay: control_delay_element  generic map(name => " 69_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(29), ack => convTransposeA_CP_4083_elements(69), clk => clk, reset =>reset);
    -- CP-element group 70:  transition  output  delay-element  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	29 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/$exit
      -- CP-element group 70: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/$exit
      -- CP-element group 70: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1513_konst_delay_trans
      -- CP-element group 70: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_req
      -- 
    phi_stmt_1509_req_5069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1509_req_5069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(70), ack => phi_stmt_1509_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(70) is a control-delay.
    cp_element_70_delay: control_delay_element  generic map(name => " 70_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(29), ack => convTransposeA_CP_4083_elements(70), clk => clk, reset =>reset);
    -- CP-element group 71:  join  transition  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	79 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_1364/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(69) & convTransposeA_CP_4083_elements(70);
      gj_convTransposeA_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	66 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Sample/ra
      -- 
    ra_5089_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_0, ack => convTransposeA_CP_4083_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	66 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/Update/ca
      -- 
    ca_5094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1508_inst_ack_1, ack => convTransposeA_CP_4083_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	78 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/$exit
      -- CP-element group 74: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/$exit
      -- CP-element group 74: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_sources/type_cast_1508/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1502/phi_stmt_1502_req
      -- 
    phi_stmt_1502_req_5095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1502_req_5095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(74), ack => phi_stmt_1502_req_1); -- 
    convTransposeA_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(72) & convTransposeA_CP_4083_elements(73);
      gj_convTransposeA_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	66 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Sample/ra
      -- 
    ra_5112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_0, ack => convTransposeA_CP_4083_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	66 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/Update/ca
      -- 
    ca_5117_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1515_inst_ack_1, ack => convTransposeA_CP_4083_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/$exit
      -- CP-element group 77: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/$exit
      -- CP-element group 77: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_sources/type_cast_1515/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_1509/phi_stmt_1509_req
      -- 
    phi_stmt_1509_req_5118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1509_req_5118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(77), ack => phi_stmt_1509_req_1); -- 
    convTransposeA_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(75) & convTransposeA_CP_4083_elements(76);
      gj_convTransposeA_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  join  transition  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	74 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1364/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeA_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(74) & convTransposeA_CP_4083_elements(77);
      gj_convTransposeA_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  merge  fork  transition  place  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	71 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1364/merge_stmt_1501_PhiReqMerge
      -- CP-element group 79: 	 branch_block_stmt_1364/merge_stmt_1501_PhiAck/$entry
      -- 
    convTransposeA_CP_4083_elements(79) <= OrReduce(convTransposeA_CP_4083_elements(71) & convTransposeA_CP_4083_elements(78));
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1364/merge_stmt_1501_PhiAck/phi_stmt_1502_ack
      -- 
    phi_stmt_1502_ack_5123_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1502_ack_0, ack => convTransposeA_CP_4083_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_1364/merge_stmt_1501_PhiAck/phi_stmt_1509_ack
      -- 
    phi_stmt_1509_ack_5124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1509_ack_0, ack => convTransposeA_CP_4083_elements(81)); -- 
    -- CP-element group 82:  join  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	30 
    -- CP-element group 82: 	31 
    -- CP-element group 82: 	32 
    -- CP-element group 82: 	33 
    -- CP-element group 82:  members (16) 
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1364/merge_stmt_1501__exit__
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629__entry__
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/$entry
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Sample/rr
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_update_start_
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1526_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Update/cr
      -- CP-element group 82: 	 branch_block_stmt_1364/assign_stmt_1522_to_assign_stmt_1629/type_cast_1521_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_1364/merge_stmt_1501_PhiAck/$exit
      -- 
    rr_4676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1521_inst_req_0); -- 
    cr_4695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1526_inst_req_1); -- 
    rr_4690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1526_inst_req_0); -- 
    cr_4681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(82), ack => type_cast_1521_inst_req_1); -- 
    convTransposeA_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(80) & convTransposeA_CP_4083_elements(81);
      gj_convTransposeA_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	57 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Sample/ra
      -- 
    ra_5144_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_0, ack => convTransposeA_CP_4083_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	57 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/Update/ca
      -- 
    ca_5149_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1638_inst_ack_1, ack => convTransposeA_CP_4083_elements(84)); -- 
    -- CP-element group 85:  join  transition  output  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (6) 
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/$exit
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$exit
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/$exit
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1638/SplitProtocol/$exit
      -- CP-element group 85: 	 branch_block_stmt_1364/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_req
      -- 
    phi_stmt_1632_req_5150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1632_req_5150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(85), ack => phi_stmt_1632_req_1); -- 
    convTransposeA_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeA_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeA_CP_4083_elements(83) & convTransposeA_CP_4083_elements(84);
      gj_convTransposeA_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeA_CP_4083_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  transition  output  delay-element  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (5) 
      -- CP-element group 86: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 86: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/$exit
      -- CP-element group 86: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/$exit
      -- CP-element group 86: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_sources/type_cast_1636_konst_delay_trans
      -- CP-element group 86: 	 branch_block_stmt_1364/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_1632/phi_stmt_1632_req
      -- 
    phi_stmt_1632_req_5161_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1632_req_5161_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(86), ack => phi_stmt_1632_req_0); -- 
    -- Element group convTransposeA_CP_4083_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => convTransposeA_CP_4083_elements(34), ack => convTransposeA_CP_4083_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  merge  transition  place  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_1364/merge_stmt_1631_PhiReqMerge
      -- CP-element group 87: 	 branch_block_stmt_1364/merge_stmt_1631_PhiAck/$entry
      -- 
    convTransposeA_CP_4083_elements(87) <= OrReduce(convTransposeA_CP_4083_elements(85) & convTransposeA_CP_4083_elements(86));
    -- CP-element group 88:  fork  transition  place  input  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	42 
    -- CP-element group 88: 	44 
    -- CP-element group 88: 	46 
    -- CP-element group 88: 	48 
    -- CP-element group 88: 	50 
    -- CP-element group 88: 	53 
    -- CP-element group 88: 	54 
    -- CP-element group 88: 	55 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	36 
    -- CP-element group 88: 	38 
    -- CP-element group 88: 	40 
    -- CP-element group 88:  members (45) 
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1690_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1716_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/merge_stmt_1631__exit__
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738__entry__
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1679_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1710_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/array_obj_ref_1685_final_index_sum_regn_update_start
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1648_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1686_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/addr_of_1717_complete/req
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/word_0/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/ptr_deref_1720_Update/word_access_complete/word_0/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1364/assign_stmt_1645_to_assign_stmt_1738/type_cast_1726_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1364/merge_stmt_1631_PhiAck/$exit
      -- CP-element group 88: 	 branch_block_stmt_1364/merge_stmt_1631_PhiAck/phi_stmt_1632_ack
      -- 
    phi_stmt_1632_ack_5166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1632_ack_0, ack => convTransposeA_CP_4083_elements(88)); -- 
    cr_4817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => ptr_deref_1690_load_0_req_1); -- 
    cr_4726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1679_inst_req_1); -- 
    cr_4836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1710_inst_req_1); -- 
    req_4867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => array_obj_ref_1716_index_offset_req_1); -- 
    req_4757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => array_obj_ref_1685_index_offset_req_1); -- 
    cr_4712_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4712_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1648_inst_req_1); -- 
    rr_4707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1648_inst_req_0); -- 
    req_4772_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4772_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => addr_of_1686_final_reg_req_1); -- 
    req_4882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_4882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => addr_of_1717_final_reg_req_1); -- 
    cr_4932_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4932_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => ptr_deref_1720_store_0_req_1); -- 
    rr_4941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_4941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1726_inst_req_0); -- 
    cr_4946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_4946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeA_CP_4083_elements(88), ack => type_cast_1726_inst_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_1591_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1612_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1672_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_1704_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1420_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1420_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom52_1715_resized : std_logic_vector(13 downto 0);
    signal R_idxprom52_1715_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_1684_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_1684_scaled : std_logic_vector(13 downto 0);
    signal add16_1552 : std_logic_vector(31 downto 0);
    signal add27_1567 : std_logic_vector(31 downto 0);
    signal add42_1624 : std_logic_vector(31 downto 0);
    signal add44_1659 : std_logic_vector(31 downto 0);
    signal add57_1733 : std_logic_vector(31 downto 0);
    signal add8_1654 : std_logic_vector(31 downto 0);
    signal add_1537 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1685_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1685_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1685_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1685_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1685_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1685_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1716_root_address : std_logic_vector(13 downto 0);
    signal arrayidx53_1718 : std_logic_vector(31 downto 0);
    signal arrayidx_1687 : std_logic_vector(31 downto 0);
    signal call_1367 : std_logic_vector(15 downto 0);
    signal cmp68_1769 : std_logic_vector(0 downto 0);
    signal cmp77_1795 : std_logic_vector(0 downto 0);
    signal cmp_1738 : std_logic_vector(0 downto 0);
    signal conv13_1406 : std_logic_vector(31 downto 0);
    signal conv18_1425 : std_logic_vector(31 downto 0);
    signal conv24_1439 : std_logic_vector(31 downto 0);
    signal conv37_1593 : std_logic_vector(31 downto 0);
    signal conv3_1522 : std_logic_vector(31 downto 0);
    signal conv40_1614 : std_logic_vector(31 downto 0);
    signal conv56_1727 : std_logic_vector(31 downto 0);
    signal conv66_1764 : std_logic_vector(31 downto 0);
    signal conv6_1527 : std_logic_vector(31 downto 0);
    signal conv74_1790 : std_logic_vector(31 downto 0);
    signal conv90_1649 : std_logic_vector(31 downto 0);
    signal div76_1499 : std_logic_vector(31 downto 0);
    signal div_1481 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1489 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1376 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1388 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1398 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1414 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1431 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1447 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1459 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1471 : std_logic_vector(31 downto 0);
    signal idxprom52_1711 : std_logic_vector(63 downto 0);
    signal idxprom_1680 : std_logic_vector(63 downto 0);
    signal inc72_1773 : std_logic_vector(15 downto 0);
    signal inc72x_xinput_dim0x_x2_1778 : std_logic_vector(15 downto 0);
    signal inc_1759 : std_logic_vector(15 downto 0);
    signal indvar_1632 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_1751 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1509 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1502 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_1785 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_1645 : std_logic_vector(15 downto 0);
    signal mul14_1547 : std_logic_vector(31 downto 0);
    signal mul25_1562 : std_logic_vector(31 downto 0);
    signal mul41_1619 : std_logic_vector(31 downto 0);
    signal mul43_1629 : std_logic_vector(31 downto 0);
    signal mul7_1542 : std_logic_vector(31 downto 0);
    signal mul_1532 : std_logic_vector(31 downto 0);
    signal ptr_deref_1379_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1379_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1379_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1379_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1379_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1391_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1391_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1391_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1391_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1391_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1401_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1401_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1401_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1401_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1401_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1417_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1417_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1417_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1417_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1417_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1434_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1434_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1434_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1434_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1434_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1450_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1450_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1450_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1450_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1450_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1462_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1462_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1462_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1462_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1462_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1474_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1474_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1474_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1474_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1474_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1492_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1492_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1492_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1492_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1492_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1690_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1690_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1690_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1720_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1720_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1720_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext91_1605 : std_logic_vector(31 downto 0);
    signal sext93_1665 : std_logic_vector(31 downto 0);
    signal sext94_1697 : std_logic_vector(31 downto 0);
    signal sext_1584 : std_logic_vector(31 downto 0);
    signal shr51_1706 : std_logic_vector(31 downto 0);
    signal shr_1674 : std_logic_vector(31 downto 0);
    signal sub19_1599 : std_logic_vector(31 downto 0);
    signal sub30_1572 : std_logic_vector(31 downto 0);
    signal sub31_1578 : std_logic_vector(31 downto 0);
    signal sub_1557 : std_logic_vector(31 downto 0);
    signal tmp12_1402 : std_logic_vector(15 downto 0);
    signal tmp15_1418 : std_logic_vector(31 downto 0);
    signal tmp17_1421 : std_logic_vector(15 downto 0);
    signal tmp1_1380 : std_logic_vector(31 downto 0);
    signal tmp23_1435 : std_logic_vector(15 downto 0);
    signal tmp26_1451 : std_logic_vector(31 downto 0);
    signal tmp35_1463 : std_logic_vector(31 downto 0);
    signal tmp38_1475 : std_logic_vector(31 downto 0);
    signal tmp48_1691 : std_logic_vector(63 downto 0);
    signal tmp4_1392 : std_logic_vector(31 downto 0);
    signal tmp75_1493 : std_logic_vector(31 downto 0);
    signal type_cast_1479_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1497_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1506_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1508_wire : std_logic_vector(15 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1515_wire : std_logic_vector(15 downto 0);
    signal type_cast_1520_wire : std_logic_vector(31 downto 0);
    signal type_cast_1525_wire : std_logic_vector(31 downto 0);
    signal type_cast_1576_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1582_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1587_wire : std_logic_vector(31 downto 0);
    signal type_cast_1590_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1603_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1608_wire : std_logic_vector(31 downto 0);
    signal type_cast_1611_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1636_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1638_wire : std_logic_vector(15 downto 0);
    signal type_cast_1643_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1663_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1668_wire : std_logic_vector(31 downto 0);
    signal type_cast_1671_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1678_wire : std_logic_vector(63 downto 0);
    signal type_cast_1695_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1700_wire : std_logic_vector(31 downto 0);
    signal type_cast_1703_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1709_wire : std_logic_vector(63 downto 0);
    signal type_cast_1725_wire : std_logic_vector(31 downto 0);
    signal type_cast_1731_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1749_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1757_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1762_wire : std_logic_vector(31 downto 0);
    signal type_cast_1782_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1788_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1420_word_address_0 <= "0";
    array_obj_ref_1685_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1685_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1685_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1685_resized_base_address <= "00000000000000";
    array_obj_ref_1716_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1716_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1716_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1716_resized_base_address <= "00000000000000";
    iNsTr_10_1489 <= "00000000000000000000000000000010";
    iNsTr_2_1376 <= "00000000000000000000000000000100";
    iNsTr_3_1388 <= "00000000000000000000000000000011";
    iNsTr_4_1398 <= "00000000000000000000000000000000";
    iNsTr_5_1414 <= "00000000000000000000000000000011";
    iNsTr_6_1431 <= "00000000000000000000000000000001";
    iNsTr_7_1447 <= "00000000000000000000000000000100";
    iNsTr_8_1459 <= "00000000000000000000000000000100";
    iNsTr_9_1471 <= "00000000000000000000000000000011";
    ptr_deref_1379_word_offset_0 <= "0000000";
    ptr_deref_1391_word_offset_0 <= "0000000";
    ptr_deref_1401_word_offset_0 <= "0";
    ptr_deref_1417_word_offset_0 <= "0000000";
    ptr_deref_1434_word_offset_0 <= "0";
    ptr_deref_1450_word_offset_0 <= "0000000";
    ptr_deref_1462_word_offset_0 <= "0000000";
    ptr_deref_1474_word_offset_0 <= "0000000";
    ptr_deref_1492_word_offset_0 <= "0000000";
    ptr_deref_1690_word_offset_0 <= "00000000000000";
    ptr_deref_1720_word_offset_0 <= "00000000000000";
    type_cast_1479_wire_constant <= "00000000000000000000000000000001";
    type_cast_1497_wire_constant <= "00000000000000000000000000000001";
    type_cast_1506_wire_constant <= "0000000000000000";
    type_cast_1513_wire_constant <= "0000000000000000";
    type_cast_1576_wire_constant <= "00000000000000000000000000010000";
    type_cast_1582_wire_constant <= "11111111111111110000000000000000";
    type_cast_1590_wire_constant <= "00000000000000000000000000010000";
    type_cast_1597_wire_constant <= "00000000000000000000000000010000";
    type_cast_1603_wire_constant <= "11111111111111110000000000000000";
    type_cast_1611_wire_constant <= "00000000000000000000000000010000";
    type_cast_1636_wire_constant <= "0000000000000000";
    type_cast_1643_wire_constant <= "0000000000000100";
    type_cast_1663_wire_constant <= "00000000000000000000000000010000";
    type_cast_1671_wire_constant <= "00000000000000000000000000010010";
    type_cast_1695_wire_constant <= "00000000000000000000000000010000";
    type_cast_1703_wire_constant <= "00000000000000000000000000010010";
    type_cast_1731_wire_constant <= "00000000000000000000000000000100";
    type_cast_1749_wire_constant <= "0000000000000001";
    type_cast_1757_wire_constant <= "0000000000000001";
    type_cast_1782_wire_constant <= "0000000000000000";
    phi_stmt_1502: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1506_wire_constant & type_cast_1508_wire;
      req <= phi_stmt_1502_req_0 & phi_stmt_1502_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1502",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1502_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1502,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1502
    phi_stmt_1509: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1513_wire_constant & type_cast_1515_wire;
      req <= phi_stmt_1509_req_0 & phi_stmt_1509_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1509",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1509_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1509,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1509
    phi_stmt_1632: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1636_wire_constant & type_cast_1638_wire;
      req <= phi_stmt_1632_req_0 & phi_stmt_1632_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1632",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1632_ack_0,
          idata => idata,
          odata => indvar_1632,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1632
    -- flow-through select operator MUX_1784_inst
    input_dim1x_x2_1785 <= type_cast_1782_wire_constant when (cmp68_1769(0) /=  '0') else inc_1759;
    addr_of_1686_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1686_final_reg_req_0;
      addr_of_1686_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1686_final_reg_req_1;
      addr_of_1686_final_reg_ack_1<= rack(0);
      addr_of_1686_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1686_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1685_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1717_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1717_final_reg_req_0;
      addr_of_1717_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1717_final_reg_req_1;
      addr_of_1717_final_reg_ack_1<= rack(0);
      addr_of_1717_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1717_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1716_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx53_1718,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1405_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1405_inst_req_0;
      type_cast_1405_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1405_inst_req_1;
      type_cast_1405_inst_ack_1<= rack(0);
      type_cast_1405_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1405_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp12_1402,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_1406,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1424_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1424_inst_req_0;
      type_cast_1424_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1424_inst_req_1;
      type_cast_1424_inst_ack_1<= rack(0);
      type_cast_1424_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1424_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp17_1421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv18_1425,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1438_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1438_inst_req_0;
      type_cast_1438_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1438_inst_req_1;
      type_cast_1438_inst_ack_1<= rack(0);
      type_cast_1438_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1438_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp23_1435,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv24_1439,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1508_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1508_inst_req_0;
      type_cast_1508_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1508_inst_req_1;
      type_cast_1508_inst_ack_1<= rack(0);
      type_cast_1508_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1508_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_1785,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1508_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1515_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1515_inst_req_0;
      type_cast_1515_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1515_inst_req_1;
      type_cast_1515_inst_ack_1<= rack(0);
      type_cast_1515_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1515_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc72x_xinput_dim0x_x2_1778,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1515_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1521_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1521_inst_req_0;
      type_cast_1521_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1521_inst_req_1;
      type_cast_1521_inst_ack_1<= rack(0);
      type_cast_1521_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1521_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1520_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv3_1522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1526_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1526_inst_req_0;
      type_cast_1526_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1526_inst_req_1;
      type_cast_1526_inst_ack_1<= rack(0);
      type_cast_1526_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1526_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1525_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv6_1527,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1587_inst
    process(sext_1584) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_1584(31 downto 0);
      type_cast_1587_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1592_inst
    process(ASHR_i32_i32_1591_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1591_wire(31 downto 0);
      conv37_1593 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1608_inst
    process(sext91_1605) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext91_1605(31 downto 0);
      type_cast_1608_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1613_inst
    process(ASHR_i32_i32_1612_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1612_wire(31 downto 0);
      conv40_1614 <= tmp_var; -- 
    end process;
    type_cast_1638_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1638_inst_req_0;
      type_cast_1638_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1638_inst_req_1;
      type_cast_1638_inst_ack_1<= rack(0);
      type_cast_1638_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1638_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1751,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1638_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1648_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1648_inst_req_0;
      type_cast_1648_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1648_inst_req_1;
      type_cast_1648_inst_ack_1<= rack(0);
      type_cast_1648_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1648_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_1645,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_1649,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1668_inst
    process(sext93_1665) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext93_1665(31 downto 0);
      type_cast_1668_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1673_inst
    process(ASHR_i32_i32_1672_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1672_wire(31 downto 0);
      shr_1674 <= tmp_var; -- 
    end process;
    type_cast_1679_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1679_inst_req_0;
      type_cast_1679_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1679_inst_req_1;
      type_cast_1679_inst_ack_1<= rack(0);
      type_cast_1679_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1679_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1678_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_1680,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1700_inst
    process(sext94_1697) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext94_1697(31 downto 0);
      type_cast_1700_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1705_inst
    process(ASHR_i32_i32_1704_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_1704_wire(31 downto 0);
      shr51_1706 <= tmp_var; -- 
    end process;
    type_cast_1710_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1710_inst_req_0;
      type_cast_1710_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1710_inst_req_1;
      type_cast_1710_inst_ack_1<= rack(0);
      type_cast_1710_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1710_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1709_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom52_1711,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1726_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1726_inst_req_0;
      type_cast_1726_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1726_inst_req_1;
      type_cast_1726_inst_ack_1<= rack(0);
      type_cast_1726_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1726_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1725_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv56_1727,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1763_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1763_inst_req_0;
      type_cast_1763_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1763_inst_req_1;
      type_cast_1763_inst_ack_1<= rack(0);
      type_cast_1763_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1763_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1762_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_1764,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1772_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1772_inst_req_0;
      type_cast_1772_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1772_inst_req_1;
      type_cast_1772_inst_ack_1<= rack(0);
      type_cast_1772_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1772_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp68_1769,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc72_1773,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1789_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1789_inst_req_0;
      type_cast_1789_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1789_inst_req_1;
      type_cast_1789_inst_ack_1<= rack(0);
      type_cast_1789_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1789_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1788_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_1790,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1420_gather_scatter
    process(LOAD_padding_1420_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1420_data_0;
      ov(15 downto 0) := iv;
      tmp17_1421 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1685_index_1_rename
    process(R_idxprom_1684_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_1684_resized;
      ov(13 downto 0) := iv;
      R_idxprom_1684_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1685_index_1_resize
    process(idxprom_1680) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_1680;
      ov := iv(13 downto 0);
      R_idxprom_1684_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1685_root_address_inst
    process(array_obj_ref_1685_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1685_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1685_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1716_index_1_rename
    process(R_idxprom52_1715_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom52_1715_resized;
      ov(13 downto 0) := iv;
      R_idxprom52_1715_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1716_index_1_resize
    process(idxprom52_1711) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom52_1711;
      ov := iv(13 downto 0);
      R_idxprom52_1715_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1716_root_address_inst
    process(array_obj_ref_1716_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1716_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1716_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1379_addr_0
    process(ptr_deref_1379_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1379_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1379_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1379_base_resize
    process(iNsTr_2_1376) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1376;
      ov := iv(6 downto 0);
      ptr_deref_1379_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1379_gather_scatter
    process(ptr_deref_1379_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1379_data_0;
      ov(31 downto 0) := iv;
      tmp1_1380 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1379_root_address_inst
    process(ptr_deref_1379_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1379_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1379_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1391_addr_0
    process(ptr_deref_1391_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1391_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1391_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1391_base_resize
    process(iNsTr_3_1388) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1388;
      ov := iv(6 downto 0);
      ptr_deref_1391_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1391_gather_scatter
    process(ptr_deref_1391_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1391_data_0;
      ov(31 downto 0) := iv;
      tmp4_1392 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1391_root_address_inst
    process(ptr_deref_1391_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1391_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1391_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1401_addr_0
    process(ptr_deref_1401_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1401_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1401_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1401_base_resize
    process(iNsTr_4_1398) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1398;
      ov := iv(0 downto 0);
      ptr_deref_1401_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1401_gather_scatter
    process(ptr_deref_1401_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1401_data_0;
      ov(15 downto 0) := iv;
      tmp12_1402 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1401_root_address_inst
    process(ptr_deref_1401_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1401_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1401_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1417_addr_0
    process(ptr_deref_1417_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1417_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1417_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1417_base_resize
    process(iNsTr_5_1414) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1414;
      ov := iv(6 downto 0);
      ptr_deref_1417_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1417_gather_scatter
    process(ptr_deref_1417_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1417_data_0;
      ov(31 downto 0) := iv;
      tmp15_1418 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1417_root_address_inst
    process(ptr_deref_1417_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1417_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1417_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1434_addr_0
    process(ptr_deref_1434_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1434_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1434_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1434_base_resize
    process(iNsTr_6_1431) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1431;
      ov := iv(0 downto 0);
      ptr_deref_1434_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1434_gather_scatter
    process(ptr_deref_1434_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1434_data_0;
      ov(15 downto 0) := iv;
      tmp23_1435 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1434_root_address_inst
    process(ptr_deref_1434_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1434_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1434_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1450_addr_0
    process(ptr_deref_1450_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1450_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1450_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1450_base_resize
    process(iNsTr_7_1447) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1447;
      ov := iv(6 downto 0);
      ptr_deref_1450_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1450_gather_scatter
    process(ptr_deref_1450_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1450_data_0;
      ov(31 downto 0) := iv;
      tmp26_1451 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1450_root_address_inst
    process(ptr_deref_1450_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1450_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1450_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_addr_0
    process(ptr_deref_1462_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1462_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1462_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_base_resize
    process(iNsTr_8_1459) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1459;
      ov := iv(6 downto 0);
      ptr_deref_1462_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_gather_scatter
    process(ptr_deref_1462_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1462_data_0;
      ov(31 downto 0) := iv;
      tmp35_1463 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1462_root_address_inst
    process(ptr_deref_1462_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1462_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1462_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_addr_0
    process(ptr_deref_1474_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1474_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1474_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_base_resize
    process(iNsTr_9_1471) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1471;
      ov := iv(6 downto 0);
      ptr_deref_1474_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_gather_scatter
    process(ptr_deref_1474_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1474_data_0;
      ov(31 downto 0) := iv;
      tmp38_1475 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1474_root_address_inst
    process(ptr_deref_1474_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1474_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1474_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1492_addr_0
    process(ptr_deref_1492_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1492_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1492_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1492_base_resize
    process(iNsTr_10_1489) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1489;
      ov := iv(6 downto 0);
      ptr_deref_1492_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1492_gather_scatter
    process(ptr_deref_1492_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1492_data_0;
      ov(31 downto 0) := iv;
      tmp75_1493 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1492_root_address_inst
    process(ptr_deref_1492_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1492_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1492_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_addr_0
    process(ptr_deref_1690_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1690_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1690_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_base_resize
    process(arrayidx_1687) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1687;
      ov := iv(13 downto 0);
      ptr_deref_1690_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_gather_scatter
    process(ptr_deref_1690_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1690_data_0;
      ov(63 downto 0) := iv;
      tmp48_1691 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1690_root_address_inst
    process(ptr_deref_1690_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1690_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1690_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_addr_0
    process(ptr_deref_1720_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1720_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_base_resize
    process(arrayidx53_1718) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx53_1718;
      ov := iv(13 downto 0);
      ptr_deref_1720_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_gather_scatter
    process(tmp48_1691) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp48_1691;
      ov(63 downto 0) := iv;
      ptr_deref_1720_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1720_root_address_inst
    process(ptr_deref_1720_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1720_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1720_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1739_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_1738;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1739_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1739_branch_req_0,
          ack0 => if_stmt_1739_branch_ack_0,
          ack1 => if_stmt_1739_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1796_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_1795;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1796_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1796_branch_req_0,
          ack0 => if_stmt_1796_branch_ack_0,
          ack1 => if_stmt_1796_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_1750_inst
    process(indvar_1632) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1632, type_cast_1749_wire_constant, tmp_var);
      indvarx_xnext_1751 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1758_inst
    process(input_dim1x_x1x_xph_1502) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1502, type_cast_1757_wire_constant, tmp_var);
      inc_1759 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_1777_inst
    process(inc72_1773, input_dim0x_x2x_xph_1509) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc72_1773, input_dim0x_x2x_xph_1509, tmp_var);
      inc72x_xinput_dim0x_x2_1778 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1536_inst
    process(mul_1532, conv3_1522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1532, conv3_1522, tmp_var);
      add_1537 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1551_inst
    process(mul14_1547, tmp15_1418) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul14_1547, tmp15_1418, tmp_var);
      add16_1552 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1566_inst
    process(mul25_1562, tmp26_1451) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul25_1562, tmp26_1451, tmp_var);
      add27_1567 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1583_inst
    process(sub31_1578) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub31_1578, type_cast_1582_wire_constant, tmp_var);
      sext_1584 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1604_inst
    process(sub19_1599) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub19_1599, type_cast_1603_wire_constant, tmp_var);
      sext91_1605 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1623_inst
    process(conv37_1593, mul41_1619) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv37_1593, mul41_1619, tmp_var);
      add42_1624 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1653_inst
    process(mul7_1542, conv90_1649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul7_1542, conv90_1649, tmp_var);
      add8_1654 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1658_inst
    process(mul43_1629, conv90_1649) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul43_1629, conv90_1649, tmp_var);
      add44_1659 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1732_inst
    process(conv56_1727) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv56_1727, type_cast_1731_wire_constant, tmp_var);
      add57_1733 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1591_inst
    process(type_cast_1587_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1587_wire, type_cast_1590_wire_constant, tmp_var);
      ASHR_i32_i32_1591_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1612_inst
    process(type_cast_1608_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1608_wire, type_cast_1611_wire_constant, tmp_var);
      ASHR_i32_i32_1612_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1672_inst
    process(type_cast_1668_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1668_wire, type_cast_1671_wire_constant, tmp_var);
      ASHR_i32_i32_1672_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_1704_inst
    process(type_cast_1700_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_1700_wire, type_cast_1703_wire_constant, tmp_var);
      ASHR_i32_i32_1704_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1768_inst
    process(conv66_1764, div_1481) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv66_1764, div_1481, tmp_var);
      cmp68_1769 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1794_inst
    process(conv74_1790, div76_1499) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv74_1790, div76_1499, tmp_var);
      cmp77_1795 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1480_inst
    process(tmp4_1392) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp4_1392, type_cast_1479_wire_constant, tmp_var);
      div_1481 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1498_inst
    process(tmp75_1493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp75_1493, type_cast_1497_wire_constant, tmp_var);
      div76_1499 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_1644_inst
    process(indvar_1632) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_1632, type_cast_1643_wire_constant, tmp_var);
      input_dim2x_x1_1645 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1531_inst
    process(tmp4_1392, conv6_1527) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp4_1392, conv6_1527, tmp_var);
      mul_1532 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1541_inst
    process(add_1537, tmp1_1380) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1537, tmp1_1380, tmp_var);
      mul7_1542 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1546_inst
    process(conv13_1406, conv6_1527) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv13_1406, conv6_1527, tmp_var);
      mul14_1547 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1561_inst
    process(conv24_1439, conv3_1522) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv24_1439, conv3_1522, tmp_var);
      mul25_1562 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1618_inst
    process(tmp38_1475, conv40_1614) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp38_1475, conv40_1614, tmp_var);
      mul41_1619 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1628_inst
    process(add42_1624, tmp35_1463) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add42_1624, tmp35_1463, tmp_var);
      mul43_1629 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1577_inst
    process(sub30_1572) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub30_1572, type_cast_1576_wire_constant, tmp_var);
      sub31_1578 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1598_inst
    process(sub_1557) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_1557, type_cast_1597_wire_constant, tmp_var);
      sub19_1599 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1664_inst
    process(add8_1654) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add8_1654, type_cast_1663_wire_constant, tmp_var);
      sext93_1665 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_1696_inst
    process(add44_1659) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add44_1659, type_cast_1695_wire_constant, tmp_var);
      sext94_1697 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1556_inst
    process(add16_1552, conv18_1425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add16_1552, conv18_1425, tmp_var);
      sub_1557 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1571_inst
    process(add27_1567, conv18_1425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add27_1567, conv18_1425, tmp_var);
      sub30_1572 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_1737_inst
    process(add57_1733, tmp1_1380) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add57_1733, tmp1_1380, tmp_var);
      cmp_1738 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_1685_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_1684_scaled;
      array_obj_ref_1685_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1685_index_offset_req_0;
      array_obj_ref_1685_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1685_index_offset_req_1;
      array_obj_ref_1685_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_1716_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom52_1715_scaled;
      array_obj_ref_1716_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1716_index_offset_req_0;
      array_obj_ref_1716_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1716_index_offset_req_1;
      array_obj_ref_1716_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_1520_inst
    process(input_dim1x_x1x_xph_1502) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1502, tmp_var);
      type_cast_1520_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1525_inst
    process(input_dim0x_x2x_xph_1509) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1509, tmp_var);
      type_cast_1525_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1678_inst
    process(shr_1674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_1674, tmp_var);
      type_cast_1678_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1709_inst
    process(shr51_1706) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr51_1706, tmp_var);
      type_cast_1709_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1725_inst
    process(input_dim2x_x1_1645) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_1645, tmp_var);
      type_cast_1725_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1762_inst
    process(inc_1759) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_1759, tmp_var);
      type_cast_1762_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1788_inst
    process(inc72x_xinput_dim0x_x2_1778) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc72x_xinput_dim0x_x2_1778, tmp_var);
      type_cast_1788_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1420_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1420_load_0_req_0;
      LOAD_padding_1420_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1420_load_0_req_1;
      LOAD_padding_1420_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1420_word_address_0;
      LOAD_padding_1420_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1379_load_0 ptr_deref_1391_load_0 ptr_deref_1492_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1379_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1391_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1492_load_0_req_0;
      ptr_deref_1379_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1391_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1492_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1379_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1391_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1492_load_0_req_1;
      ptr_deref_1379_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1391_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1492_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1379_word_address_0 & ptr_deref_1391_word_address_0 & ptr_deref_1492_word_address_0;
      ptr_deref_1379_data_0 <= data_out(95 downto 64);
      ptr_deref_1391_data_0 <= data_out(63 downto 32);
      ptr_deref_1492_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1401_load_0 ptr_deref_1434_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1401_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1434_load_0_req_0;
      ptr_deref_1401_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1434_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1401_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1434_load_0_req_1;
      ptr_deref_1401_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1434_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1401_word_address_0 & ptr_deref_1434_word_address_0;
      ptr_deref_1401_data_0 <= data_out(31 downto 16);
      ptr_deref_1434_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1417_load_0 ptr_deref_1450_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1417_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1450_load_0_req_0;
      ptr_deref_1417_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1450_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1417_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1450_load_0_req_1;
      ptr_deref_1417_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1450_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1417_word_address_0 & ptr_deref_1450_word_address_0;
      ptr_deref_1417_data_0 <= data_out(63 downto 32);
      ptr_deref_1450_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1462_load_0 ptr_deref_1474_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1462_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1474_load_0_req_0;
      ptr_deref_1462_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1474_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1462_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1474_load_0_req_1;
      ptr_deref_1462_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1474_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1462_word_address_0 & ptr_deref_1474_word_address_0;
      ptr_deref_1462_data_0 <= data_out(63 downto 32);
      ptr_deref_1474_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_1690_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1690_load_0_req_0;
      ptr_deref_1690_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1690_load_0_req_1;
      ptr_deref_1690_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1690_word_address_0;
      ptr_deref_1690_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_1720_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1720_store_0_req_0;
      ptr_deref_1720_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1720_store_0_req_1;
      ptr_deref_1720_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1720_word_address_0;
      data_in <= ptr_deref_1720_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block0_start_1366_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block0_start_1366_inst_req_0;
      RPIPE_Block0_start_1366_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block0_start_1366_inst_req_1;
      RPIPE_Block0_start_1366_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1367 <= data_out(15 downto 0);
      Block0_start_read_0_gI: SplitGuardInterface generic map(name => "Block0_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block0_start_read_0: InputPortRevised -- 
        generic map ( name => "Block0_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block0_start_pipe_read_req(0),
          oack => Block0_start_pipe_read_ack(0),
          odata => Block0_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block0_done_1804_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block0_done_1804_inst_req_0;
      WPIPE_Block0_done_1804_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block0_done_1804_inst_req_1;
      WPIPE_Block0_done_1804_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1367;
      Block0_done_write_0_gI: SplitGuardInterface generic map(name => "Block0_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block0_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block0_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block0_done_pipe_write_req(0),
          oack => Block0_done_pipe_write_ack(0),
          odata => Block0_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeA_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeB is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeB;
architecture convTransposeB_arch of convTransposeB is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeB_CP_5207_start: Boolean;
  signal convTransposeB_CP_5207_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_1875_load_0_ack_1 : boolean;
  signal LOAD_padding_1878_load_0_req_1 : boolean;
  signal type_cast_1882_inst_ack_1 : boolean;
  signal type_cast_1882_inst_req_1 : boolean;
  signal LOAD_padding_1878_load_0_ack_1 : boolean;
  signal ptr_deref_1875_load_0_req_1 : boolean;
  signal type_cast_1882_inst_ack_0 : boolean;
  signal ptr_deref_1908_load_0_req_1 : boolean;
  signal ptr_deref_1908_load_0_ack_1 : boolean;
  signal type_cast_1896_inst_req_0 : boolean;
  signal type_cast_1896_inst_ack_0 : boolean;
  signal ptr_deref_1892_load_0_req_0 : boolean;
  signal ptr_deref_1892_load_0_ack_0 : boolean;
  signal ptr_deref_1892_load_0_req_1 : boolean;
  signal LOAD_padding_1878_load_0_req_0 : boolean;
  signal ptr_deref_1892_load_0_ack_1 : boolean;
  signal LOAD_padding_1878_load_0_ack_0 : boolean;
  signal ptr_deref_1908_load_0_req_0 : boolean;
  signal ptr_deref_1908_load_0_ack_0 : boolean;
  signal type_cast_1896_inst_req_1 : boolean;
  signal type_cast_1896_inst_ack_1 : boolean;
  signal type_cast_1882_inst_req_0 : boolean;
  signal ptr_deref_1875_load_0_req_0 : boolean;
  signal ptr_deref_1875_load_0_ack_0 : boolean;
  signal ptr_deref_1920_load_0_req_0 : boolean;
  signal ptr_deref_1920_load_0_ack_0 : boolean;
  signal RPIPE_Block1_start_1814_inst_req_0 : boolean;
  signal RPIPE_Block1_start_1814_inst_ack_0 : boolean;
  signal RPIPE_Block1_start_1814_inst_req_1 : boolean;
  signal RPIPE_Block1_start_1814_inst_ack_1 : boolean;
  signal ptr_deref_1827_load_0_req_0 : boolean;
  signal ptr_deref_1827_load_0_ack_0 : boolean;
  signal ptr_deref_1827_load_0_req_1 : boolean;
  signal ptr_deref_1827_load_0_ack_1 : boolean;
  signal type_cast_1837_inst_req_0 : boolean;
  signal type_cast_1837_inst_ack_0 : boolean;
  signal type_cast_1837_inst_req_1 : boolean;
  signal type_cast_1837_inst_ack_1 : boolean;
  signal ptr_deref_1849_load_0_req_0 : boolean;
  signal ptr_deref_1849_load_0_ack_0 : boolean;
  signal ptr_deref_1849_load_0_req_1 : boolean;
  signal ptr_deref_1849_load_0_ack_1 : boolean;
  signal ptr_deref_1859_load_0_req_0 : boolean;
  signal ptr_deref_1859_load_0_ack_0 : boolean;
  signal ptr_deref_1859_load_0_req_1 : boolean;
  signal ptr_deref_1859_load_0_ack_1 : boolean;
  signal type_cast_1863_inst_req_0 : boolean;
  signal type_cast_1863_inst_ack_0 : boolean;
  signal type_cast_1863_inst_req_1 : boolean;
  signal type_cast_1863_inst_ack_1 : boolean;
  signal ptr_deref_1920_load_0_req_1 : boolean;
  signal ptr_deref_1920_load_0_ack_1 : boolean;
  signal ptr_deref_1932_load_0_req_0 : boolean;
  signal ptr_deref_1932_load_0_ack_0 : boolean;
  signal ptr_deref_1932_load_0_req_1 : boolean;
  signal ptr_deref_1932_load_0_ack_1 : boolean;
  signal ptr_deref_1944_load_0_req_0 : boolean;
  signal ptr_deref_1944_load_0_ack_0 : boolean;
  signal ptr_deref_1944_load_0_req_1 : boolean;
  signal ptr_deref_1944_load_0_ack_1 : boolean;
  signal type_cast_1971_inst_req_0 : boolean;
  signal type_cast_1971_inst_ack_0 : boolean;
  signal type_cast_1971_inst_req_1 : boolean;
  signal type_cast_1971_inst_ack_1 : boolean;
  signal type_cast_1976_inst_req_0 : boolean;
  signal type_cast_1976_inst_ack_0 : boolean;
  signal type_cast_1976_inst_req_1 : boolean;
  signal type_cast_1976_inst_ack_1 : boolean;
  signal type_cast_2098_inst_req_0 : boolean;
  signal type_cast_2098_inst_ack_0 : boolean;
  signal type_cast_2098_inst_req_1 : boolean;
  signal type_cast_2098_inst_ack_1 : boolean;
  signal type_cast_2128_inst_req_0 : boolean;
  signal type_cast_2128_inst_ack_0 : boolean;
  signal type_cast_2128_inst_req_1 : boolean;
  signal type_cast_2128_inst_ack_1 : boolean;
  signal array_obj_ref_2134_index_offset_req_0 : boolean;
  signal array_obj_ref_2134_index_offset_ack_0 : boolean;
  signal array_obj_ref_2134_index_offset_req_1 : boolean;
  signal array_obj_ref_2134_index_offset_ack_1 : boolean;
  signal addr_of_2135_final_reg_req_0 : boolean;
  signal addr_of_2135_final_reg_ack_0 : boolean;
  signal addr_of_2135_final_reg_req_1 : boolean;
  signal addr_of_2135_final_reg_ack_1 : boolean;
  signal ptr_deref_2139_load_0_req_0 : boolean;
  signal ptr_deref_2139_load_0_ack_0 : boolean;
  signal ptr_deref_2139_load_0_req_1 : boolean;
  signal ptr_deref_2139_load_0_ack_1 : boolean;
  signal type_cast_2159_inst_req_0 : boolean;
  signal type_cast_2159_inst_ack_0 : boolean;
  signal type_cast_2159_inst_req_1 : boolean;
  signal type_cast_2159_inst_ack_1 : boolean;
  signal array_obj_ref_2165_index_offset_req_0 : boolean;
  signal array_obj_ref_2165_index_offset_ack_0 : boolean;
  signal array_obj_ref_2165_index_offset_req_1 : boolean;
  signal array_obj_ref_2165_index_offset_ack_1 : boolean;
  signal addr_of_2166_final_reg_req_0 : boolean;
  signal addr_of_2166_final_reg_ack_0 : boolean;
  signal addr_of_2166_final_reg_req_1 : boolean;
  signal addr_of_2166_final_reg_ack_1 : boolean;
  signal ptr_deref_2169_store_0_req_0 : boolean;
  signal ptr_deref_2169_store_0_ack_0 : boolean;
  signal ptr_deref_2169_store_0_req_1 : boolean;
  signal ptr_deref_2169_store_0_ack_1 : boolean;
  signal type_cast_2175_inst_req_0 : boolean;
  signal type_cast_2175_inst_ack_0 : boolean;
  signal type_cast_2175_inst_req_1 : boolean;
  signal type_cast_2175_inst_ack_1 : boolean;
  signal if_stmt_2188_branch_req_0 : boolean;
  signal if_stmt_2188_branch_ack_1 : boolean;
  signal if_stmt_2188_branch_ack_0 : boolean;
  signal type_cast_2212_inst_req_0 : boolean;
  signal type_cast_2212_inst_ack_0 : boolean;
  signal type_cast_2212_inst_req_1 : boolean;
  signal type_cast_2212_inst_ack_1 : boolean;
  signal if_stmt_2219_branch_req_0 : boolean;
  signal if_stmt_2219_branch_ack_1 : boolean;
  signal if_stmt_2219_branch_ack_0 : boolean;
  signal type_cast_2240_inst_req_0 : boolean;
  signal type_cast_2240_inst_ack_0 : boolean;
  signal type_cast_2240_inst_req_1 : boolean;
  signal type_cast_2240_inst_ack_1 : boolean;
  signal type_cast_2260_inst_req_0 : boolean;
  signal type_cast_2260_inst_ack_0 : boolean;
  signal type_cast_2260_inst_req_1 : boolean;
  signal type_cast_2260_inst_ack_1 : boolean;
  signal if_stmt_2267_branch_req_0 : boolean;
  signal if_stmt_2267_branch_ack_1 : boolean;
  signal if_stmt_2267_branch_ack_0 : boolean;
  signal WPIPE_Block1_done_2275_inst_req_0 : boolean;
  signal WPIPE_Block1_done_2275_inst_ack_0 : boolean;
  signal WPIPE_Block1_done_2275_inst_req_1 : boolean;
  signal WPIPE_Block1_done_2275_inst_ack_1 : boolean;
  signal phi_stmt_1960_req_0 : boolean;
  signal type_cast_1957_inst_req_0 : boolean;
  signal type_cast_1957_inst_ack_0 : boolean;
  signal type_cast_1957_inst_req_1 : boolean;
  signal type_cast_1957_inst_ack_1 : boolean;
  signal phi_stmt_1954_req_0 : boolean;
  signal type_cast_1966_inst_req_0 : boolean;
  signal type_cast_1966_inst_ack_0 : boolean;
  signal type_cast_1966_inst_req_1 : boolean;
  signal type_cast_1966_inst_ack_1 : boolean;
  signal phi_stmt_1960_req_1 : boolean;
  signal type_cast_1959_inst_req_0 : boolean;
  signal type_cast_1959_inst_ack_0 : boolean;
  signal type_cast_1959_inst_req_1 : boolean;
  signal type_cast_1959_inst_ack_1 : boolean;
  signal phi_stmt_1954_req_1 : boolean;
  signal phi_stmt_1954_ack_0 : boolean;
  signal phi_stmt_1960_ack_0 : boolean;
  signal type_cast_2085_inst_req_0 : boolean;
  signal type_cast_2085_inst_ack_0 : boolean;
  signal type_cast_2085_inst_req_1 : boolean;
  signal type_cast_2085_inst_ack_1 : boolean;
  signal phi_stmt_2082_req_0 : boolean;
  signal phi_stmt_2082_req_1 : boolean;
  signal phi_stmt_2082_ack_0 : boolean;
  signal type_cast_2249_inst_req_0 : boolean;
  signal type_cast_2249_inst_ack_0 : boolean;
  signal type_cast_2249_inst_req_1 : boolean;
  signal type_cast_2249_inst_ack_1 : boolean;
  signal phi_stmt_2244_req_1 : boolean;
  signal type_cast_2255_inst_req_0 : boolean;
  signal type_cast_2255_inst_ack_0 : boolean;
  signal type_cast_2255_inst_req_1 : boolean;
  signal type_cast_2255_inst_ack_1 : boolean;
  signal phi_stmt_2250_req_1 : boolean;
  signal type_cast_2247_inst_req_0 : boolean;
  signal type_cast_2247_inst_ack_0 : boolean;
  signal type_cast_2247_inst_req_1 : boolean;
  signal type_cast_2247_inst_ack_1 : boolean;
  signal phi_stmt_2244_req_0 : boolean;
  signal type_cast_2253_inst_req_0 : boolean;
  signal type_cast_2253_inst_ack_0 : boolean;
  signal type_cast_2253_inst_req_1 : boolean;
  signal type_cast_2253_inst_ack_1 : boolean;
  signal phi_stmt_2250_req_0 : boolean;
  signal phi_stmt_2244_ack_0 : boolean;
  signal phi_stmt_2250_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeB_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeB_CP_5207_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeB_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeB_CP_5207_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeB_CP_5207: Block -- control-path 
    signal convTransposeB_CP_5207_elements: BooleanArray(112 downto 0);
    -- 
  begin -- 
    convTransposeB_CP_5207_elements(0) <= convTransposeB_CP_5207_start;
    convTransposeB_CP_5207_symbol <= convTransposeB_CP_5207_elements(72);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1812/$entry
      -- CP-element group 0: 	 branch_block_stmt_1812/branch_block_stmt_1812__entry__
      -- CP-element group 0: 	 branch_block_stmt_1812/assign_stmt_1815__entry__
      -- CP-element group 0: 	 branch_block_stmt_1812/assign_stmt_1815/$entry
      -- CP-element group 0: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Sample/rr
      -- 
    rr_5265_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5265_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(0), ack => RPIPE_Block1_start_1814_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_update_start_
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Update/cr
      -- 
    ra_5266_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1814_inst_ack_0, ack => convTransposeB_CP_5207_elements(1)); -- 
    cr_5270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(1), ack => RPIPE_Block1_start_1814_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1815__exit__
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951__entry__
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1815/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1815/RPIPE_Block1_start_1814_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_update_start_
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/word_0/cr
      -- 
    ca_5271_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block1_start_1814_inst_ack_1, ack => convTransposeB_CP_5207_elements(2)); -- 
    cr_5529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => LOAD_padding_1878_load_0_req_1); -- 
    cr_5548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1882_inst_req_1); -- 
    cr_5496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1875_load_0_req_1); -- 
    cr_5657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1908_load_0_req_1); -- 
    rr_5582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1892_load_0_req_0); -- 
    cr_5593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1892_load_0_req_1); -- 
    rr_5518_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5518_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => LOAD_padding_1878_load_0_req_0); -- 
    rr_5646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1908_load_0_req_0); -- 
    cr_5612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1896_inst_req_1); -- 
    rr_5485_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5485_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1875_load_0_req_0); -- 
    rr_5696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1920_load_0_req_0); -- 
    rr_5307_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5307_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1827_load_0_req_0); -- 
    cr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1827_load_0_req_1); -- 
    cr_5337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1837_inst_req_1); -- 
    rr_5371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1849_load_0_req_0); -- 
    cr_5382_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5382_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1849_load_0_req_1); -- 
    rr_5421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1859_load_0_req_0); -- 
    cr_5432_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5432_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1859_load_0_req_1); -- 
    cr_5451_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5451_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => type_cast_1863_inst_req_1); -- 
    cr_5707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1920_load_0_req_1); -- 
    rr_5746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1932_load_0_req_0); -- 
    cr_5757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1932_load_0_req_1); -- 
    rr_5796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1944_load_0_req_0); -- 
    cr_5807_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5807_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(2), ack => ptr_deref_1944_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Sample/word_access_start/word_0/ra
      -- 
    ra_5308_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1827_load_0_ack_0, ack => convTransposeB_CP_5207_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/ptr_deref_1827_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/ptr_deref_1827_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/ptr_deref_1827_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1827_Update/ptr_deref_1827_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Sample/rr
      -- 
    ca_5319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1827_load_0_ack_1, ack => convTransposeB_CP_5207_elements(4)); -- 
    rr_5332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(4), ack => type_cast_1837_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Sample/ra
      -- 
    ra_5333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_0, ack => convTransposeB_CP_5207_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1837_Update/ca
      -- 
    ca_5338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1837_inst_ack_1, ack => convTransposeB_CP_5207_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Sample/word_access_start/word_0/ra
      -- 
    ra_5372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1849_load_0_ack_0, ack => convTransposeB_CP_5207_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/ptr_deref_1849_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/ptr_deref_1849_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/ptr_deref_1849_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1849_Update/ptr_deref_1849_Merge/merge_ack
      -- 
    ca_5383_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1849_load_0_ack_1, ack => convTransposeB_CP_5207_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/$exit
      -- CP-element group 9: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Sample/word_access_start/word_0/ra
      -- 
    ra_5422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1859_load_0_ack_0, ack => convTransposeB_CP_5207_elements(9)); -- 
    -- CP-element group 10:  transition  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10:  members (12) 
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/ptr_deref_1859_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/ptr_deref_1859_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/ptr_deref_1859_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1859_Update/ptr_deref_1859_Merge/merge_ack
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_sample_start_
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Sample/rr
      -- 
    ca_5433_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1859_load_0_ack_1, ack => convTransposeB_CP_5207_elements(10)); -- 
    rr_5446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(10), ack => type_cast_1863_inst_req_0); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Sample/ra
      -- 
    ra_5447_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_0, ack => convTransposeB_CP_5207_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	31 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1863_Update/ca
      -- 
    ca_5452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1863_inst_ack_1, ack => convTransposeB_CP_5207_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Sample/word_access_start/word_0/ra
      -- CP-element group 13: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_sample_completed_
      -- 
    ra_5486_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1875_load_0_ack_0, ack => convTransposeB_CP_5207_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (9) 
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/ptr_deref_1875_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/ptr_deref_1875_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/ptr_deref_1875_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_Update/ptr_deref_1875_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1875_update_completed_
      -- 
    ca_5497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1875_load_0_ack_1, ack => convTransposeB_CP_5207_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/word_access_start/word_0/ra
      -- CP-element group 15: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Sample/$exit
      -- 
    ra_5519_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1878_load_0_ack_0, ack => convTransposeB_CP_5207_elements(15)); -- 
    -- CP-element group 16:  transition  input  output  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (12) 
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_sample_start_
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Sample/$entry
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/LOAD_padding_1878_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Sample/rr
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/LOAD_padding_1878_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/LOAD_padding_1878_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/LOAD_padding_1878_Update/LOAD_padding_1878_Merge/merge_ack
      -- 
    ca_5530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_1878_load_0_ack_1, ack => convTransposeB_CP_5207_elements(16)); -- 
    rr_5543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(16), ack => type_cast_1882_inst_req_0); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Sample/ra
      -- CP-element group 17: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Sample/$exit
      -- 
    ra_5544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_0, ack => convTransposeB_CP_5207_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	31 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Update/ca
      -- CP-element group 18: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1882_Update/$exit
      -- 
    ca_5549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1882_inst_ack_1, ack => convTransposeB_CP_5207_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Sample/word_access_start/word_0/ra
      -- 
    ra_5583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1892_load_0_ack_0, ack => convTransposeB_CP_5207_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/ptr_deref_1892_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/ptr_deref_1892_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/ptr_deref_1892_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/ptr_deref_1892_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1892_Update/$exit
      -- 
    ca_5594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1892_load_0_ack_1, ack => convTransposeB_CP_5207_elements(20)); -- 
    rr_5607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(20), ack => type_cast_1896_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_sample_completed_
      -- 
    ra_5608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_0, ack => convTransposeB_CP_5207_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/type_cast_1896_update_completed_
      -- 
    ca_5613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_1, ack => convTransposeB_CP_5207_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_sample_completed_
      -- 
    ra_5647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1908_load_0_ack_0, ack => convTransposeB_CP_5207_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (9) 
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/ptr_deref_1908_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/ptr_deref_1908_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/ptr_deref_1908_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_Update/ptr_deref_1908_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1908_update_completed_
      -- 
    ca_5658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1908_load_0_ack_1, ack => convTransposeB_CP_5207_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Sample/word_access_start/word_0/ra
      -- 
    ra_5697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1920_load_0_ack_0, ack => convTransposeB_CP_5207_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/ptr_deref_1920_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/ptr_deref_1920_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/ptr_deref_1920_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1920_Update/ptr_deref_1920_Merge/merge_ack
      -- 
    ca_5708_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1920_load_0_ack_1, ack => convTransposeB_CP_5207_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Sample/word_access_start/word_0/ra
      -- 
    ra_5747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1932_load_0_ack_0, ack => convTransposeB_CP_5207_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/ptr_deref_1932_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/ptr_deref_1932_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/ptr_deref_1932_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1932_Update/ptr_deref_1932_Merge/merge_ack
      -- 
    ca_5758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1932_load_0_ack_1, ack => convTransposeB_CP_5207_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Sample/word_access_start/word_0/ra
      -- 
    ra_5797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1944_load_0_ack_0, ack => convTransposeB_CP_5207_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/ptr_deref_1944_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/ptr_deref_1944_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/ptr_deref_1944_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/ptr_deref_1944_Update/ptr_deref_1944_Merge/merge_ack
      -- 
    ca_5808_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1944_load_0_ack_1, ack => convTransposeB_CP_5207_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	12 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	18 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	8 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	73 
    -- CP-element group 31: 	74 
    -- CP-element group 31: 	75 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951__exit__
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_1812/assign_stmt_1824_to_assign_stmt_1951/$exit
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/cr
      -- 
    rr_6250_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6250_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(31), ack => type_cast_1957_inst_req_0); -- 
    cr_6255_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6255_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(31), ack => type_cast_1957_inst_req_1); -- 
    convTransposeB_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(12) & convTransposeB_CP_5207_elements(22) & convTransposeB_CP_5207_elements(24) & convTransposeB_CP_5207_elements(26) & convTransposeB_CP_5207_elements(28) & convTransposeB_CP_5207_elements(30) & convTransposeB_CP_5207_elements(18) & convTransposeB_CP_5207_elements(14) & convTransposeB_CP_5207_elements(6) & convTransposeB_CP_5207_elements(8);
      gj_convTransposeB_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	88 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Sample/ra
      -- 
    ra_5825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_0, ack => convTransposeB_CP_5207_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	88 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Update/ca
      -- 
    ca_5830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1971_inst_ack_1, ack => convTransposeB_CP_5207_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	88 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Sample/ra
      -- 
    ra_5839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_0, ack => convTransposeB_CP_5207_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	88 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Update/ca
      -- 
    ca_5844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1976_inst_ack_1, ack => convTransposeB_CP_5207_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	92 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079__exit__
      -- CP-element group 36: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/$exit
      -- CP-element group 36: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/$entry
      -- CP-element group 36: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/$entry
      -- 
    convTransposeB_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(35) & convTransposeB_CP_5207_elements(33);
      gj_convTransposeB_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	94 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Sample/ra
      -- 
    ra_5856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2098_inst_ack_0, ack => convTransposeB_CP_5207_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	94 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Sample/rr
      -- 
    ca_5861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2098_inst_ack_1, ack => convTransposeB_CP_5207_elements(38)); -- 
    rr_5869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(38), ack => type_cast_2128_inst_req_0); -- 
    rr_5979_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5979_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(38), ack => type_cast_2159_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Sample/ra
      -- 
    ra_5870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_0, ack => convTransposeB_CP_5207_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	94 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Sample/req
      -- 
    ca_5875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2128_inst_ack_1, ack => convTransposeB_CP_5207_elements(40)); -- 
    req_5900_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5900_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(40), ack => array_obj_ref_2134_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Sample/ack
      -- 
    ack_5901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2134_index_offset_ack_0, ack => convTransposeB_CP_5207_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	94 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_request/req
      -- 
    ack_5906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2134_index_offset_ack_1, ack => convTransposeB_CP_5207_elements(42)); -- 
    req_5915_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5915_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(42), ack => addr_of_2135_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_request/ack
      -- 
    ack_5916_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2135_final_reg_ack_0, ack => convTransposeB_CP_5207_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	94 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/word_0/rr
      -- 
    ack_5921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2135_final_reg_ack_1, ack => convTransposeB_CP_5207_elements(44)); -- 
    rr_5954_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5954_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(44), ack => ptr_deref_2139_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Sample/word_access_start/word_0/ra
      -- 
    ra_5955_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2139_load_0_ack_0, ack => convTransposeB_CP_5207_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	94 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/ptr_deref_2139_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/ptr_deref_2139_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/ptr_deref_2139_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/ptr_deref_2139_Merge/merge_ack
      -- 
    ca_5966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2139_load_0_ack_1, ack => convTransposeB_CP_5207_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Sample/ra
      -- 
    ra_5980_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2159_inst_ack_0, ack => convTransposeB_CP_5207_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	94 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Sample/req
      -- 
    ca_5985_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2159_inst_ack_1, ack => convTransposeB_CP_5207_elements(48)); -- 
    req_6010_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6010_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(48), ack => array_obj_ref_2165_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Sample/ack
      -- 
    ack_6011_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2165_index_offset_ack_0, ack => convTransposeB_CP_5207_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	94 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_base_plus_offset/sum_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_request/req
      -- 
    ack_6016_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2165_index_offset_ack_1, ack => convTransposeB_CP_5207_elements(50)); -- 
    req_6025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(50), ack => addr_of_2166_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_request/ack
      -- 
    ack_6026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2166_final_reg_ack_0, ack => convTransposeB_CP_5207_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	94 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_word_addrgen/root_register_ack
      -- 
    ack_6031_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2166_final_reg_ack_1, ack => convTransposeB_CP_5207_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	46 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/ptr_deref_2169_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/ptr_deref_2169_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/ptr_deref_2169_Split/split_req
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/ptr_deref_2169_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/word_0/rr
      -- 
    rr_6069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(53), ack => ptr_deref_2169_store_0_req_0); -- 
    convTransposeB_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(46) & convTransposeB_CP_5207_elements(52);
      gj_convTransposeB_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/$exit
      -- CP-element group 54: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Sample/word_access_start/word_0/ra
      -- 
    ra_6070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_store_0_ack_0, ack => convTransposeB_CP_5207_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	94 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/$exit
      -- CP-element group 55: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/word_0/ca
      -- 
    ca_6081_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2169_store_0_ack_1, ack => convTransposeB_CP_5207_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	94 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Sample/ra
      -- 
    ra_6090_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2175_inst_ack_0, ack => convTransposeB_CP_5207_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	94 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Update/ca
      -- 
    ca_6095_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2175_inst_ack_1, ack => convTransposeB_CP_5207_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	55 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187__exit__
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188__entry__
      -- CP-element group 58: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/$exit
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_1812/R_cmp_2189_place
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_1812/if_stmt_2188_else_link/$entry
      -- 
    branch_req_6103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(58), ack => if_stmt_2188_branch_req_0); -- 
    convTransposeB_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(41) & convTransposeB_CP_5207_elements(49) & convTransposeB_CP_5207_elements(57) & convTransposeB_CP_5207_elements(55);
      gj_convTransposeB_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	89 
    -- CP-element group 59: 	90 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_1812/merge_stmt_2194__exit__
      -- CP-element group 59: 	 branch_block_stmt_1812/assign_stmt_2200__entry__
      -- CP-element group 59: 	 branch_block_stmt_1812/assign_stmt_2200__exit__
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_1812/if_stmt_2188_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1812/if_stmt_2188_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1812/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_1812/assign_stmt_2200/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/assign_stmt_2200/$exit
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_1812/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_1812/merge_stmt_2194_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_1812/merge_stmt_2194_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_1812/merge_stmt_2194_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_1812/merge_stmt_2194_PhiAck/dummy
      -- 
    if_choice_transition_6108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2188_branch_ack_1, ack => convTransposeB_CP_5207_elements(59)); -- 
    rr_6331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(59), ack => type_cast_2085_inst_req_0); -- 
    cr_6336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(59), ack => type_cast_2085_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	61 
    -- CP-element group 60:  members (18) 
      -- CP-element group 60: 	 branch_block_stmt_1812/merge_stmt_2202__exit__
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218__entry__
      -- CP-element group 60: 	 branch_block_stmt_1812/if_stmt_2188_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_1812/if_stmt_2188_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_1812/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/$entry
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_update_start_
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_1812/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_1812/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1812/merge_stmt_2202_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_1812/merge_stmt_2202_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_1812/merge_stmt_2202_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_1812/merge_stmt_2202_PhiAck/dummy
      -- 
    else_choice_transition_6112_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2188_branch_ack_0, ack => convTransposeB_CP_5207_elements(60)); -- 
    rr_6128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(60), ack => type_cast_2212_inst_req_0); -- 
    cr_6133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(60), ack => type_cast_2212_inst_req_1); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Sample/ra
      -- 
    ra_6129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2212_inst_ack_0, ack => convTransposeB_CP_5207_elements(61)); -- 
    -- CP-element group 62:  branch  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (13) 
      -- CP-element group 62: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218__exit__
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219__entry__
      -- CP-element group 62: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/$exit
      -- CP-element group 62: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1812/assign_stmt_2208_to_assign_stmt_2218/type_cast_2212_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_dead_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_eval_test/$entry
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_eval_test/$exit
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_eval_test/branch_req
      -- CP-element group 62: 	 branch_block_stmt_1812/R_cmp77_2220_place
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_if_link/$entry
      -- CP-element group 62: 	 branch_block_stmt_1812/if_stmt_2219_else_link/$entry
      -- 
    ca_6134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2212_inst_ack_1, ack => convTransposeB_CP_5207_elements(62)); -- 
    branch_req_6142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(62), ack => if_stmt_2219_branch_req_0); -- 
    -- CP-element group 63:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	66 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (18) 
      -- CP-element group 63: 	 branch_block_stmt_1812/merge_stmt_2225__exit__
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241__entry__
      -- CP-element group 63: 	 branch_block_stmt_1812/if_stmt_2219_if_link/$exit
      -- CP-element group 63: 	 branch_block_stmt_1812/if_stmt_2219_if_link/if_choice_transition
      -- CP-element group 63: 	 branch_block_stmt_1812/ifx_xelse_ifx_xthen79
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/$entry
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Sample/rr
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Update/cr
      -- CP-element group 63: 	 branch_block_stmt_1812/ifx_xelse_ifx_xthen79_PhiReq/$entry
      -- CP-element group 63: 	 branch_block_stmt_1812/ifx_xelse_ifx_xthen79_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1812/merge_stmt_2225_PhiReqMerge
      -- CP-element group 63: 	 branch_block_stmt_1812/merge_stmt_2225_PhiAck/$entry
      -- CP-element group 63: 	 branch_block_stmt_1812/merge_stmt_2225_PhiAck/$exit
      -- CP-element group 63: 	 branch_block_stmt_1812/merge_stmt_2225_PhiAck/dummy
      -- 
    if_choice_transition_6147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2219_branch_ack_1, ack => convTransposeB_CP_5207_elements(63)); -- 
    rr_6164_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6164_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(63), ack => type_cast_2240_inst_req_0); -- 
    cr_6169_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6169_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(63), ack => type_cast_2240_inst_req_1); -- 
    -- CP-element group 64:  fork  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	95 
    -- CP-element group 64: 	96 
    -- CP-element group 64: 	99 
    -- CP-element group 64: 	98 
    -- CP-element group 64:  members (20) 
      -- CP-element group 64: 	 branch_block_stmt_1812/if_stmt_2219_else_link/$exit
      -- CP-element group 64: 	 branch_block_stmt_1812/if_stmt_2219_else_link/else_choice_transition
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Update/cr
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Update/$entry
      -- CP-element group 64: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2219_branch_ack_0, ack => convTransposeB_CP_5207_elements(64)); -- 
    rr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2249_inst_req_0); -- 
    cr_6410_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6410_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2249_inst_req_1); -- 
    rr_6428_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6428_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2255_inst_req_0); -- 
    cr_6433_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6433_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(64), ack => type_cast_2255_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Sample/ra
      -- 
    ra_6165_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2240_inst_ack_0, ack => convTransposeB_CP_5207_elements(65)); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	63 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	106 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66: 	105 
    -- CP-element group 66:  members (23) 
      -- CP-element group 66: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241__exit__
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/$exit
      -- CP-element group 66: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_1812/assign_stmt_2231_to_assign_stmt_2241/type_cast_2240_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Update/cr
      -- 
    ca_6170_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2240_inst_ack_1, ack => convTransposeB_CP_5207_elements(66)); -- 
    rr_6454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2247_inst_req_0); -- 
    cr_6459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2247_inst_req_1); -- 
    rr_6477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2253_inst_req_0); -- 
    cr_6482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(66), ack => type_cast_2253_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	112 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Sample/ra
      -- 
    ra_6182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_0, ack => convTransposeB_CP_5207_elements(67)); -- 
    -- CP-element group 68:  branch  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	112 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (13) 
      -- CP-element group 68: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266__exit__
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267__entry__
      -- CP-element group 68: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/$exit
      -- CP-element group 68: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_dead_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_eval_test/$entry
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_eval_test/$exit
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_eval_test/branch_req
      -- CP-element group 68: 	 branch_block_stmt_1812/R_cmp89_2268_place
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_if_link/$entry
      -- CP-element group 68: 	 branch_block_stmt_1812/if_stmt_2267_else_link/$entry
      -- 
    ca_6187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2260_inst_ack_1, ack => convTransposeB_CP_5207_elements(68)); -- 
    branch_req_6195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_6195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(68), ack => if_stmt_2267_branch_req_0); -- 
    -- CP-element group 69:  merge  transition  place  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (15) 
      -- CP-element group 69: 	 branch_block_stmt_1812/merge_stmt_2273__exit__
      -- CP-element group 69: 	 branch_block_stmt_1812/assign_stmt_2277__entry__
      -- CP-element group 69: 	 branch_block_stmt_1812/if_stmt_2267_if_link/$exit
      -- CP-element group 69: 	 branch_block_stmt_1812/if_stmt_2267_if_link/if_choice_transition
      -- CP-element group 69: 	 branch_block_stmt_1812/ifx_xend_whilex_xend
      -- CP-element group 69: 	 branch_block_stmt_1812/assign_stmt_2277/$entry
      -- CP-element group 69: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Sample/$entry
      -- CP-element group 69: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Sample/req
      -- CP-element group 69: 	 branch_block_stmt_1812/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 69: 	 branch_block_stmt_1812/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 69: 	 branch_block_stmt_1812/merge_stmt_2273_PhiReqMerge
      -- CP-element group 69: 	 branch_block_stmt_1812/merge_stmt_2273_PhiAck/$entry
      -- CP-element group 69: 	 branch_block_stmt_1812/merge_stmt_2273_PhiAck/$exit
      -- CP-element group 69: 	 branch_block_stmt_1812/merge_stmt_2273_PhiAck/dummy
      -- 
    if_choice_transition_6200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2267_branch_ack_1, ack => convTransposeB_CP_5207_elements(69)); -- 
    req_6217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(69), ack => WPIPE_Block1_done_2275_inst_req_0); -- 
    -- CP-element group 70:  fork  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	78 
    -- CP-element group 70: 	79 
    -- CP-element group 70: 	81 
    -- CP-element group 70: 	82 
    -- CP-element group 70:  members (20) 
      -- CP-element group 70: 	 branch_block_stmt_1812/if_stmt_2267_else_link/$exit
      -- CP-element group 70: 	 branch_block_stmt_1812/if_stmt_2267_else_link/else_choice_transition
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Update/cr
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Sample/rr
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Update/$entry
      -- CP-element group 70: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Update/cr
      -- 
    else_choice_transition_6204_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2267_branch_ack_0, ack => convTransposeB_CP_5207_elements(70)); -- 
    rr_6276_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6276_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1966_inst_req_0); -- 
    cr_6281_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6281_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1966_inst_req_1); -- 
    rr_6299_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6299_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1959_inst_req_0); -- 
    cr_6304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(70), ack => type_cast_1959_inst_req_1); -- 
    -- CP-element group 71:  transition  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Update/req
      -- 
    ack_6218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2275_inst_ack_0, ack => convTransposeB_CP_5207_elements(71)); -- 
    req_6222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(71), ack => WPIPE_Block1_done_2275_inst_req_1); -- 
    -- CP-element group 72:  transition  place  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72:  members (16) 
      -- CP-element group 72: 	 $exit
      -- CP-element group 72: 	 branch_block_stmt_1812/$exit
      -- CP-element group 72: 	 branch_block_stmt_1812/branch_block_stmt_1812__exit__
      -- CP-element group 72: 	 branch_block_stmt_1812/assign_stmt_2277__exit__
      -- CP-element group 72: 	 branch_block_stmt_1812/return__
      -- CP-element group 72: 	 branch_block_stmt_1812/merge_stmt_2279__exit__
      -- CP-element group 72: 	 branch_block_stmt_1812/assign_stmt_2277/$exit
      -- CP-element group 72: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_1812/assign_stmt_2277/WPIPE_Block1_done_2275_Update/ack
      -- CP-element group 72: 	 branch_block_stmt_1812/return___PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_1812/return___PhiReq/$exit
      -- CP-element group 72: 	 branch_block_stmt_1812/merge_stmt_2279_PhiReqMerge
      -- CP-element group 72: 	 branch_block_stmt_1812/merge_stmt_2279_PhiAck/$entry
      -- CP-element group 72: 	 branch_block_stmt_1812/merge_stmt_2279_PhiAck/$exit
      -- CP-element group 72: 	 branch_block_stmt_1812/merge_stmt_2279_PhiAck/dummy
      -- 
    ack_6223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block1_done_2275_inst_ack_1, ack => convTransposeB_CP_5207_elements(72)); -- 
    -- CP-element group 73:  transition  output  delay-element  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	77 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/$exit
      -- CP-element group 73: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/$exit
      -- CP-element group 73: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1964_konst_delay_trans
      -- CP-element group 73: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_req
      -- 
    phi_stmt_1960_req_6234_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1960_req_6234_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(73), ack => phi_stmt_1960_req_0); -- 
    -- Element group convTransposeB_CP_5207_elements(73) is a control-delay.
    cp_element_73_delay: control_delay_element  generic map(name => " 73_delay", delay_value => 1)  port map(req => convTransposeB_CP_5207_elements(31), ack => convTransposeB_CP_5207_elements(73), clk => clk, reset =>reset);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	31 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Sample/ra
      -- 
    ra_6251_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_0, ack => convTransposeB_CP_5207_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	31 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	76 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/Update/ca
      -- 
    ca_6256_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1957_inst_ack_1, ack => convTransposeB_CP_5207_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	75 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (5) 
      -- CP-element group 76: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/$exit
      -- CP-element group 76: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$exit
      -- CP-element group 76: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/$exit
      -- CP-element group 76: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1957/SplitProtocol/$exit
      -- CP-element group 76: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_req
      -- 
    phi_stmt_1954_req_6257_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1954_req_6257_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(76), ack => phi_stmt_1954_req_0); -- 
    convTransposeB_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(74) & convTransposeB_CP_5207_elements(75);
      gj_convTransposeB_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	73 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	85 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_1812/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(73) & convTransposeB_CP_5207_elements(76);
      gj_convTransposeB_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	70 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Sample/ra
      -- 
    ra_6277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1966_inst_ack_0, ack => convTransposeB_CP_5207_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	70 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/Update/ca
      -- 
    ca_6282_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1966_inst_ack_1, ack => convTransposeB_CP_5207_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	84 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/$exit
      -- CP-element group 80: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/$exit
      -- CP-element group 80: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_sources/type_cast_1966/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1960/phi_stmt_1960_req
      -- 
    phi_stmt_1960_req_6283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1960_req_6283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(80), ack => phi_stmt_1960_req_1); -- 
    convTransposeB_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(78) & convTransposeB_CP_5207_elements(79);
      gj_convTransposeB_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	70 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Sample/ra
      -- 
    ra_6300_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_0, ack => convTransposeB_CP_5207_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	70 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/Update/ca
      -- 
    ca_6305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1959_inst_ack_1, ack => convTransposeB_CP_5207_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (5) 
      -- CP-element group 83: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/$exit
      -- CP-element group 83: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/$exit
      -- CP-element group 83: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/$exit
      -- CP-element group 83: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_sources/type_cast_1959/SplitProtocol/$exit
      -- CP-element group 83: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_1954/phi_stmt_1954_req
      -- 
    phi_stmt_1954_req_6306_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1954_req_6306_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(83), ack => phi_stmt_1954_req_1); -- 
    convTransposeB_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(81) & convTransposeB_CP_5207_elements(82);
      gj_convTransposeB_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	80 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_1812/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(80) & convTransposeB_CP_5207_elements(83);
      gj_convTransposeB_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  merge  fork  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: 	77 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_1812/merge_stmt_1953_PhiReqMerge
      -- CP-element group 85: 	 branch_block_stmt_1812/merge_stmt_1953_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(85) <= OrReduce(convTransposeB_CP_5207_elements(84) & convTransposeB_CP_5207_elements(77));
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	88 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1812/merge_stmt_1953_PhiAck/phi_stmt_1954_ack
      -- 
    phi_stmt_1954_ack_6311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1954_ack_0, ack => convTransposeB_CP_5207_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1812/merge_stmt_1953_PhiAck/phi_stmt_1960_ack
      -- 
    phi_stmt_1960_ack_6312_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1960_ack_0, ack => convTransposeB_CP_5207_elements(87)); -- 
    -- CP-element group 88:  join  fork  transition  place  output  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	86 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	34 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	32 
    -- CP-element group 88: 	33 
    -- CP-element group 88:  members (16) 
      -- CP-element group 88: 	 branch_block_stmt_1812/merge_stmt_1953__exit__
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079__entry__
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/$entry
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1971_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Sample/rr
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_1812/assign_stmt_1972_to_assign_stmt_2079/type_cast_1976_Update/cr
      -- CP-element group 88: 	 branch_block_stmt_1812/merge_stmt_1953_PhiAck/$exit
      -- 
    rr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1971_inst_req_0); -- 
    cr_5829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1971_inst_req_1); -- 
    rr_5838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1976_inst_req_0); -- 
    cr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(88), ack => type_cast_1976_inst_req_1); -- 
    convTransposeB_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(86) & convTransposeB_CP_5207_elements(87);
      gj_convTransposeB_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	59 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Sample/ra
      -- 
    ra_6332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2085_inst_ack_0, ack => convTransposeB_CP_5207_elements(89)); -- 
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	59 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (2) 
      -- CP-element group 90: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/Update/ca
      -- 
    ca_6337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2085_inst_ack_1, ack => convTransposeB_CP_5207_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2085/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1812/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_req
      -- 
    phi_stmt_2082_req_6338_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2082_req_6338_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(91), ack => phi_stmt_2082_req_0); -- 
    convTransposeB_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(89) & convTransposeB_CP_5207_elements(90);
      gj_convTransposeB_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  transition  output  delay-element  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	36 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	93 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 92: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/$exit
      -- CP-element group 92: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/$exit
      -- CP-element group 92: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_sources/type_cast_2088_konst_delay_trans
      -- CP-element group 92: 	 branch_block_stmt_1812/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2082/phi_stmt_2082_req
      -- 
    phi_stmt_2082_req_6349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2082_req_6349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(92), ack => phi_stmt_2082_req_1); -- 
    -- Element group convTransposeB_CP_5207_elements(92) is a control-delay.
    cp_element_92_delay: control_delay_element  generic map(name => " 92_delay", delay_value => 1)  port map(req => convTransposeB_CP_5207_elements(36), ack => convTransposeB_CP_5207_elements(92), clk => clk, reset =>reset);
    -- CP-element group 93:  merge  transition  place  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: 	92 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_1812/merge_stmt_2081_PhiReqMerge
      -- CP-element group 93: 	 branch_block_stmt_1812/merge_stmt_2081_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(93) <= OrReduce(convTransposeB_CP_5207_elements(91) & convTransposeB_CP_5207_elements(92));
    -- CP-element group 94:  fork  transition  place  input  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	93 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	42 
    -- CP-element group 94: 	48 
    -- CP-element group 94: 	37 
    -- CP-element group 94: 	38 
    -- CP-element group 94: 	50 
    -- CP-element group 94: 	56 
    -- CP-element group 94: 	57 
    -- CP-element group 94: 	40 
    -- CP-element group 94: 	46 
    -- CP-element group 94: 	44 
    -- CP-element group 94: 	52 
    -- CP-element group 94: 	55 
    -- CP-element group 94:  members (45) 
      -- CP-element group 94: 	 branch_block_stmt_1812/merge_stmt_2081__exit__
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187__entry__
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2098_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2128_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2134_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2135_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2139_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2159_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_update_start
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/array_obj_ref_2165_final_index_sum_regn_Update/req
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/addr_of_2166_complete/req
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/ptr_deref_2169_Update/word_access_complete/word_0/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_update_start_
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Sample/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Sample/rr
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Update/$entry
      -- CP-element group 94: 	 branch_block_stmt_1812/assign_stmt_2095_to_assign_stmt_2187/type_cast_2175_Update/cr
      -- CP-element group 94: 	 branch_block_stmt_1812/merge_stmt_2081_PhiAck/$exit
      -- CP-element group 94: 	 branch_block_stmt_1812/merge_stmt_2081_PhiAck/phi_stmt_2082_ack
      -- 
    phi_stmt_2082_ack_6354_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2082_ack_0, ack => convTransposeB_CP_5207_elements(94)); -- 
    rr_5855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_5855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2098_inst_req_0); -- 
    cr_5860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2098_inst_req_1); -- 
    cr_5874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2128_inst_req_1); -- 
    req_5905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => array_obj_ref_2134_index_offset_req_1); -- 
    req_5920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_5920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => addr_of_2135_final_reg_req_1); -- 
    cr_5965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => ptr_deref_2139_load_0_req_1); -- 
    cr_5984_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_5984_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2159_inst_req_1); -- 
    req_6015_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6015_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => array_obj_ref_2165_index_offset_req_1); -- 
    req_6030_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_6030_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => addr_of_2166_final_reg_req_1); -- 
    cr_6080_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6080_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => ptr_deref_2169_store_0_req_1); -- 
    rr_6089_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6089_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2175_inst_req_0); -- 
    cr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6094_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(94), ack => type_cast_2175_inst_req_1); -- 
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	64 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (2) 
      -- CP-element group 95: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Sample/$exit
      -- CP-element group 95: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Sample/ra
      -- 
    ra_6406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2249_inst_ack_0, ack => convTransposeB_CP_5207_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	64 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (2) 
      -- CP-element group 96: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/Update/ca
      -- 
    ca_6411_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2249_inst_ack_1, ack => convTransposeB_CP_5207_elements(96)); -- 
    -- CP-element group 97:  join  transition  output  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	101 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/$exit
      -- CP-element group 97: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/$exit
      -- CP-element group 97: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/$exit
      -- CP-element group 97: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2249/SplitProtocol/$exit
      -- CP-element group 97: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_req
      -- 
    phi_stmt_2244_req_6412_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2244_req_6412_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(97), ack => phi_stmt_2244_req_1); -- 
    convTransposeB_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeB_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(95) & convTransposeB_CP_5207_elements(96);
      gj_convTransposeB_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	64 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	100 
    -- CP-element group 98:  members (2) 
      -- CP-element group 98: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Sample/ra
      -- 
    ra_6429_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_0, ack => convTransposeB_CP_5207_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	64 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/Update/ca
      -- 
    ca_6434_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2255_inst_ack_1, ack => convTransposeB_CP_5207_elements(99)); -- 
    -- CP-element group 100:  join  transition  output  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: 	98 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (5) 
      -- CP-element group 100: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/$exit
      -- CP-element group 100: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/$exit
      -- CP-element group 100: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/$exit
      -- CP-element group 100: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2255/SplitProtocol/$exit
      -- CP-element group 100: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_req
      -- 
    phi_stmt_2250_req_6435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2250_req_6435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(100), ack => phi_stmt_2250_req_1); -- 
    convTransposeB_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(99) & convTransposeB_CP_5207_elements(98);
      gj_convTransposeB_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  join  transition  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: 	97 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	109 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_1812/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(100) & convTransposeB_CP_5207_elements(97);
      gj_convTransposeB_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Sample/ra
      -- 
    ra_6455_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_0, ack => convTransposeB_CP_5207_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/Update/ca
      -- 
    ca_6460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2247_inst_ack_1, ack => convTransposeB_CP_5207_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	108 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/$exit
      -- CP-element group 104: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/$exit
      -- CP-element group 104: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_sources/type_cast_2247/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2244/phi_stmt_2244_req
      -- 
    phi_stmt_2244_req_6461_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2244_req_6461_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(104), ack => phi_stmt_2244_req_0); -- 
    convTransposeB_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(102) & convTransposeB_CP_5207_elements(103);
      gj_convTransposeB_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	66 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	107 
    -- CP-element group 105:  members (2) 
      -- CP-element group 105: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Sample/ra
      -- 
    ra_6478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_0, ack => convTransposeB_CP_5207_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	66 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	107 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/Update/ca
      -- 
    ca_6483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2253_inst_ack_1, ack => convTransposeB_CP_5207_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	106 
    -- CP-element group 107: 	105 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (5) 
      -- CP-element group 107: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/$exit
      -- CP-element group 107: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/$exit
      -- CP-element group 107: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/$exit
      -- CP-element group 107: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_sources/type_cast_2253/SplitProtocol/$exit
      -- CP-element group 107: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/phi_stmt_2250/phi_stmt_2250_req
      -- 
    phi_stmt_2250_req_6484_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2250_req_6484_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(107), ack => phi_stmt_2250_req_0); -- 
    convTransposeB_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(106) & convTransposeB_CP_5207_elements(105);
      gj_convTransposeB_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	104 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	109 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_1812/ifx_xthen79_ifx_xend_PhiReq/$exit
      -- 
    convTransposeB_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(107) & convTransposeB_CP_5207_elements(104);
      gj_convTransposeB_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  merge  fork  transition  place  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	101 
    -- CP-element group 109: 	108 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	110 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_1812/merge_stmt_2243_PhiReqMerge
      -- CP-element group 109: 	 branch_block_stmt_1812/merge_stmt_2243_PhiAck/$entry
      -- 
    convTransposeB_CP_5207_elements(109) <= OrReduce(convTransposeB_CP_5207_elements(101) & convTransposeB_CP_5207_elements(108));
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	109 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (1) 
      -- CP-element group 110: 	 branch_block_stmt_1812/merge_stmt_2243_PhiAck/phi_stmt_2244_ack
      -- 
    phi_stmt_2244_ack_6489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2244_ack_0, ack => convTransposeB_CP_5207_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_1812/merge_stmt_2243_PhiAck/phi_stmt_2250_ack
      -- 
    phi_stmt_2250_ack_6490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2250_ack_0, ack => convTransposeB_CP_5207_elements(111)); -- 
    -- CP-element group 112:  join  fork  transition  place  output  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: 	111 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	67 
    -- CP-element group 112: 	68 
    -- CP-element group 112:  members (10) 
      -- CP-element group 112: 	 branch_block_stmt_1812/merge_stmt_2243__exit__
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266__entry__
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/$entry
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_sample_start_
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_update_start_
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Sample/$entry
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Sample/rr
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_1812/assign_stmt_2261_to_assign_stmt_2266/type_cast_2260_Update/cr
      -- CP-element group 112: 	 branch_block_stmt_1812/merge_stmt_2243_PhiAck/$exit
      -- 
    rr_6181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(112), ack => type_cast_2260_inst_req_0); -- 
    cr_6186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeB_CP_5207_elements(112), ack => type_cast_2260_inst_req_1); -- 
    convTransposeB_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeB_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeB_CP_5207_elements(110) & convTransposeB_CP_5207_elements(111);
      gj_convTransposeB_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeB_CP_5207_elements(112), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2041_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2062_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2122_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2153_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_1878_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_1878_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom61_2164_resized : std_logic_vector(13 downto 0);
    signal R_idxprom61_2164_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2133_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2133_scaled : std_logic_vector(13 downto 0);
    signal add17_2104 : std_logic_vector(31 downto 0);
    signal add25_2002 : std_logic_vector(31 downto 0);
    signal add36_2017 : std_logic_vector(31 downto 0);
    signal add51_2074 : std_logic_vector(31 downto 0);
    signal add53_2109 : std_logic_vector(31 downto 0);
    signal add66_2182 : std_logic_vector(31 downto 0);
    signal add_1987 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2134_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2134_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2134_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2134_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2134_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2134_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2165_root_address : std_logic_vector(13 downto 0);
    signal arrayidx62_2167 : std_logic_vector(31 downto 0);
    signal arrayidx_2136 : std_logic_vector(31 downto 0);
    signal call_1815 : std_logic_vector(15 downto 0);
    signal cmp77_2218 : std_logic_vector(0 downto 0);
    signal cmp89_2266 : std_logic_vector(0 downto 0);
    signal cmp_2187 : std_logic_vector(0 downto 0);
    signal conv12_1972 : std_logic_vector(31 downto 0);
    signal conv15_1977 : std_logic_vector(31 downto 0);
    signal conv22_1864 : std_logic_vector(31 downto 0);
    signal conv27_1883 : std_logic_vector(31 downto 0);
    signal conv33_1897 : std_logic_vector(31 downto 0);
    signal conv46_2043 : std_logic_vector(31 downto 0);
    signal conv49_2064 : std_logic_vector(31 downto 0);
    signal conv65_2176 : std_logic_vector(31 downto 0);
    signal conv75_2213 : std_logic_vector(31 downto 0);
    signal conv84_2241 : std_logic_vector(15 downto 0);
    signal conv86_2261 : std_logic_vector(31 downto 0);
    signal conv9102_2099 : std_logic_vector(31 downto 0);
    signal conv_1838 : std_logic_vector(15 downto 0);
    signal div83_2237 : std_logic_vector(31 downto 0);
    signal div88_1951 : std_logic_vector(31 downto 0);
    signal div_1834 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1941 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1824 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1846 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1856 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1872 : std_logic_vector(31 downto 0);
    signal iNsTr_6_1889 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1905 : std_logic_vector(31 downto 0);
    signal iNsTr_8_1917 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1929 : std_logic_vector(31 downto 0);
    signal idxprom61_2160 : std_logic_vector(63 downto 0);
    signal idxprom_2129 : std_logic_vector(63 downto 0);
    signal inc81_2231 : std_logic_vector(15 downto 0);
    signal inc_2208 : std_logic_vector(15 downto 0);
    signal indvar_2082 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2200 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_2250 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_1960 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_1954 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2244 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2095 : std_logic_vector(15 downto 0);
    signal mul16_1992 : std_logic_vector(31 downto 0);
    signal mul23_1997 : std_logic_vector(31 downto 0);
    signal mul34_2012 : std_logic_vector(31 downto 0);
    signal mul50_2069 : std_logic_vector(31 downto 0);
    signal mul52_2079 : std_logic_vector(31 downto 0);
    signal mul_1982 : std_logic_vector(31 downto 0);
    signal ptr_deref_1827_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1827_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1827_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1827_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1827_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1849_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1849_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1849_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1849_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1849_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1859_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1859_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1859_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1859_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1859_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1875_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1875_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1875_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1875_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1875_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1892_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1892_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1892_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1892_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1892_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1908_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1908_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1908_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1908_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1908_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1920_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1920_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1920_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1920_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1920_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1932_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1932_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1932_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1932_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1932_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1944_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1944_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1944_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1944_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1944_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2139_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2139_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2139_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2139_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2139_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2169_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2169_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2169_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext103_2055 : std_logic_vector(31 downto 0);
    signal sext105_2115 : std_logic_vector(31 downto 0);
    signal sext106_2146 : std_logic_vector(31 downto 0);
    signal sext_2034 : std_logic_vector(31 downto 0);
    signal shr60_2155 : std_logic_vector(31 downto 0);
    signal shr_2124 : std_logic_vector(31 downto 0);
    signal sub28_2049 : std_logic_vector(31 downto 0);
    signal sub39_2022 : std_logic_vector(31 downto 0);
    signal sub40_2028 : std_logic_vector(31 downto 0);
    signal sub_2007 : std_logic_vector(31 downto 0);
    signal tmp10_1850 : std_logic_vector(31 downto 0);
    signal tmp21_1860 : std_logic_vector(15 downto 0);
    signal tmp24_1876 : std_logic_vector(31 downto 0);
    signal tmp26_1879 : std_logic_vector(15 downto 0);
    signal tmp32_1893 : std_logic_vector(15 downto 0);
    signal tmp35_1909 : std_logic_vector(31 downto 0);
    signal tmp44_1921 : std_logic_vector(31 downto 0);
    signal tmp47_1933 : std_logic_vector(31 downto 0);
    signal tmp57_2140 : std_logic_vector(63 downto 0);
    signal tmp87_1945 : std_logic_vector(31 downto 0);
    signal tmp_1828 : std_logic_vector(31 downto 0);
    signal type_cast_1832_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1949_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1957_wire : std_logic_vector(15 downto 0);
    signal type_cast_1959_wire : std_logic_vector(15 downto 0);
    signal type_cast_1964_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1966_wire : std_logic_vector(15 downto 0);
    signal type_cast_1970_wire : std_logic_vector(31 downto 0);
    signal type_cast_1975_wire : std_logic_vector(31 downto 0);
    signal type_cast_2026_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2032_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2037_wire : std_logic_vector(31 downto 0);
    signal type_cast_2040_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2047_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2053_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2058_wire : std_logic_vector(31 downto 0);
    signal type_cast_2061_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2085_wire : std_logic_vector(15 downto 0);
    signal type_cast_2088_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2093_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2113_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2118_wire : std_logic_vector(31 downto 0);
    signal type_cast_2121_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2127_wire : std_logic_vector(63 downto 0);
    signal type_cast_2144_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2149_wire : std_logic_vector(31 downto 0);
    signal type_cast_2152_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2158_wire : std_logic_vector(63 downto 0);
    signal type_cast_2174_wire : std_logic_vector(31 downto 0);
    signal type_cast_2180_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2198_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2206_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2211_wire : std_logic_vector(31 downto 0);
    signal type_cast_2229_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2235_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2247_wire : std_logic_vector(15 downto 0);
    signal type_cast_2249_wire : std_logic_vector(15 downto 0);
    signal type_cast_2253_wire : std_logic_vector(15 downto 0);
    signal type_cast_2255_wire : std_logic_vector(15 downto 0);
    signal type_cast_2259_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_1878_word_address_0 <= "0";
    array_obj_ref_2134_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2134_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2134_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2134_resized_base_address <= "00000000000000";
    array_obj_ref_2165_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2165_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2165_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2165_resized_base_address <= "00000000000000";
    iNsTr_10_1941 <= "00000000000000000000000000000010";
    iNsTr_2_1824 <= "00000000000000000000000000000011";
    iNsTr_3_1846 <= "00000000000000000000000000000100";
    iNsTr_4_1856 <= "00000000000000000000000000000000";
    iNsTr_5_1872 <= "00000000000000000000000000000011";
    iNsTr_6_1889 <= "00000000000000000000000000000001";
    iNsTr_7_1905 <= "00000000000000000000000000000100";
    iNsTr_8_1917 <= "00000000000000000000000000000100";
    iNsTr_9_1929 <= "00000000000000000000000000000011";
    ptr_deref_1827_word_offset_0 <= "0000000";
    ptr_deref_1849_word_offset_0 <= "0000000";
    ptr_deref_1859_word_offset_0 <= "0";
    ptr_deref_1875_word_offset_0 <= "0000000";
    ptr_deref_1892_word_offset_0 <= "0";
    ptr_deref_1908_word_offset_0 <= "0000000";
    ptr_deref_1920_word_offset_0 <= "0000000";
    ptr_deref_1932_word_offset_0 <= "0000000";
    ptr_deref_1944_word_offset_0 <= "0000000";
    ptr_deref_2139_word_offset_0 <= "00000000000000";
    ptr_deref_2169_word_offset_0 <= "00000000000000";
    type_cast_1832_wire_constant <= "00000000000000000000000000000001";
    type_cast_1949_wire_constant <= "00000000000000000000000000000001";
    type_cast_1964_wire_constant <= "0000000000000000";
    type_cast_2026_wire_constant <= "00000000000000000000000000010000";
    type_cast_2032_wire_constant <= "11111111111111110000000000000000";
    type_cast_2040_wire_constant <= "00000000000000000000000000010000";
    type_cast_2047_wire_constant <= "00000000000000000000000000010000";
    type_cast_2053_wire_constant <= "11111111111111110000000000000000";
    type_cast_2061_wire_constant <= "00000000000000000000000000010000";
    type_cast_2088_wire_constant <= "0000000000000000";
    type_cast_2093_wire_constant <= "0000000000000100";
    type_cast_2113_wire_constant <= "00000000000000000000000000010000";
    type_cast_2121_wire_constant <= "00000000000000000000000000010010";
    type_cast_2144_wire_constant <= "00000000000000000000000000010000";
    type_cast_2152_wire_constant <= "00000000000000000000000000010010";
    type_cast_2180_wire_constant <= "00000000000000000000000000000100";
    type_cast_2198_wire_constant <= "0000000000000001";
    type_cast_2206_wire_constant <= "0000000000000001";
    type_cast_2229_wire_constant <= "0000000000000001";
    type_cast_2235_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1954: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1957_wire & type_cast_1959_wire;
      req <= phi_stmt_1954_req_0 & phi_stmt_1954_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1954",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1954_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_1954,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1954
    phi_stmt_1960: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1964_wire_constant & type_cast_1966_wire;
      req <= phi_stmt_1960_req_0 & phi_stmt_1960_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1960",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1960_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_1960,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1960
    phi_stmt_2082: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2085_wire & type_cast_2088_wire_constant;
      req <= phi_stmt_2082_req_0 & phi_stmt_2082_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2082",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2082_ack_0,
          idata => idata,
          odata => indvar_2082,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2082
    phi_stmt_2244: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2247_wire & type_cast_2249_wire;
      req <= phi_stmt_2244_req_0 & phi_stmt_2244_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2244",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2244_ack_0,
          idata => idata,
          odata => input_dim1x_x2_2244,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2244
    phi_stmt_2250: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2253_wire & type_cast_2255_wire;
      req <= phi_stmt_2250_req_0 & phi_stmt_2250_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2250",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2250_ack_0,
          idata => idata,
          odata => input_dim0x_x0_2250,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2250
    addr_of_2135_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2135_final_reg_req_0;
      addr_of_2135_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2135_final_reg_req_1;
      addr_of_2135_final_reg_ack_1<= rack(0);
      addr_of_2135_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2135_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2134_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2166_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2166_final_reg_req_0;
      addr_of_2166_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2166_final_reg_req_1;
      addr_of_2166_final_reg_ack_1<= rack(0);
      addr_of_2166_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2166_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2165_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx62_2167,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1837_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1837_inst_req_0;
      type_cast_1837_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1837_inst_req_1;
      type_cast_1837_inst_ack_1<= rack(0);
      type_cast_1837_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1837_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_1834,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1838,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1863_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1863_inst_req_0;
      type_cast_1863_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1863_inst_req_1;
      type_cast_1863_inst_ack_1<= rack(0);
      type_cast_1863_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1863_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp21_1860,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv22_1864,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1882_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1882_inst_req_0;
      type_cast_1882_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1882_inst_req_1;
      type_cast_1882_inst_ack_1<= rack(0);
      type_cast_1882_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1882_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp26_1879,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv27_1883,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1896_inst_req_0;
      type_cast_1896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1896_inst_req_1;
      type_cast_1896_inst_ack_1<= rack(0);
      type_cast_1896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp32_1893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv33_1897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1957_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1957_inst_req_0;
      type_cast_1957_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1957_inst_req_1;
      type_cast_1957_inst_ack_1<= rack(0);
      type_cast_1957_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1957_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_1838,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1957_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1959_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1959_inst_req_0;
      type_cast_1959_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1959_inst_req_1;
      type_cast_1959_inst_ack_1<= rack(0);
      type_cast_1959_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1959_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2244,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1959_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1966_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1966_inst_req_0;
      type_cast_1966_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1966_inst_req_1;
      type_cast_1966_inst_ack_1<= rack(0);
      type_cast_1966_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1966_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_2250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1966_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1971_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1971_inst_req_0;
      type_cast_1971_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1971_inst_req_1;
      type_cast_1971_inst_ack_1<= rack(0);
      type_cast_1971_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1971_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1970_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv12_1972,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1976_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1976_inst_req_0;
      type_cast_1976_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1976_inst_req_1;
      type_cast_1976_inst_ack_1<= rack(0);
      type_cast_1976_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1976_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_1975_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv15_1977,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2037_inst
    process(sext_2034) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2034(31 downto 0);
      type_cast_2037_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2042_inst
    process(ASHR_i32_i32_2041_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2041_wire(31 downto 0);
      conv46_2043 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2058_inst
    process(sext103_2055) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2055(31 downto 0);
      type_cast_2058_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2063_inst
    process(ASHR_i32_i32_2062_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2062_wire(31 downto 0);
      conv49_2064 <= tmp_var; -- 
    end process;
    type_cast_2085_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2085_inst_req_0;
      type_cast_2085_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2085_inst_req_1;
      type_cast_2085_inst_ack_1<= rack(0);
      type_cast_2085_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2085_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2200,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2085_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2098_inst_req_0;
      type_cast_2098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2098_inst_req_1;
      type_cast_2098_inst_ack_1<= rack(0);
      type_cast_2098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2095,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv9102_2099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2118_inst
    process(sext105_2115) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext105_2115(31 downto 0);
      type_cast_2118_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2123_inst
    process(ASHR_i32_i32_2122_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2122_wire(31 downto 0);
      shr_2124 <= tmp_var; -- 
    end process;
    type_cast_2128_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2128_inst_req_0;
      type_cast_2128_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2128_inst_req_1;
      type_cast_2128_inst_ack_1<= rack(0);
      type_cast_2128_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2128_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2127_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2129,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2149_inst
    process(sext106_2146) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2146(31 downto 0);
      type_cast_2149_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2154_inst
    process(ASHR_i32_i32_2153_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2153_wire(31 downto 0);
      shr60_2155 <= tmp_var; -- 
    end process;
    type_cast_2159_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2159_inst_req_0;
      type_cast_2159_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2159_inst_req_1;
      type_cast_2159_inst_ack_1<= rack(0);
      type_cast_2159_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2159_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2158_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom61_2160,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2175_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2175_inst_req_0;
      type_cast_2175_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2175_inst_req_1;
      type_cast_2175_inst_ack_1<= rack(0);
      type_cast_2175_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2175_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2174_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv65_2176,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2212_inst_req_0;
      type_cast_2212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2212_inst_req_1;
      type_cast_2212_inst_ack_1<= rack(0);
      type_cast_2212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2211_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv75_2213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2240_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2240_inst_req_0;
      type_cast_2240_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2240_inst_req_1;
      type_cast_2240_inst_ack_1<= rack(0);
      type_cast_2240_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2240_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div83_2237,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv84_2241,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2247_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2247_inst_req_0;
      type_cast_2247_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2247_inst_req_1;
      type_cast_2247_inst_ack_1<= rack(0);
      type_cast_2247_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2247_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv84_2241,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2247_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2249_inst_req_0;
      type_cast_2249_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2249_inst_req_1;
      type_cast_2249_inst_ack_1<= rack(0);
      type_cast_2249_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_2208,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2249_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2253_inst_req_0;
      type_cast_2253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2253_inst_req_1;
      type_cast_2253_inst_ack_1<= rack(0);
      type_cast_2253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc81_2231,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2253_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2255_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2255_inst_req_0;
      type_cast_2255_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2255_inst_req_1;
      type_cast_2255_inst_ack_1<= rack(0);
      type_cast_2255_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2255_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_1960,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2255_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2260_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2260_inst_req_0;
      type_cast_2260_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2260_inst_req_1;
      type_cast_2260_inst_ack_1<= rack(0);
      type_cast_2260_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2260_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2259_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv86_2261,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_1878_gather_scatter
    process(LOAD_padding_1878_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_1878_data_0;
      ov(15 downto 0) := iv;
      tmp26_1879 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2134_index_1_rename
    process(R_idxprom_2133_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2133_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2133_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2134_index_1_resize
    process(idxprom_2129) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2129;
      ov := iv(13 downto 0);
      R_idxprom_2133_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2134_root_address_inst
    process(array_obj_ref_2134_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2134_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2134_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2165_index_1_rename
    process(R_idxprom61_2164_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom61_2164_resized;
      ov(13 downto 0) := iv;
      R_idxprom61_2164_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2165_index_1_resize
    process(idxprom61_2160) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom61_2160;
      ov := iv(13 downto 0);
      R_idxprom61_2164_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2165_root_address_inst
    process(array_obj_ref_2165_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2165_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2165_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1827_addr_0
    process(ptr_deref_1827_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1827_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1827_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1827_base_resize
    process(iNsTr_2_1824) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1824;
      ov := iv(6 downto 0);
      ptr_deref_1827_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1827_gather_scatter
    process(ptr_deref_1827_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1827_data_0;
      ov(31 downto 0) := iv;
      tmp_1828 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1827_root_address_inst
    process(ptr_deref_1827_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1827_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1827_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1849_addr_0
    process(ptr_deref_1849_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1849_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1849_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1849_base_resize
    process(iNsTr_3_1846) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_1846;
      ov := iv(6 downto 0);
      ptr_deref_1849_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1849_gather_scatter
    process(ptr_deref_1849_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1849_data_0;
      ov(31 downto 0) := iv;
      tmp10_1850 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1849_root_address_inst
    process(ptr_deref_1849_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1849_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1849_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1859_addr_0
    process(ptr_deref_1859_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1859_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1859_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1859_base_resize
    process(iNsTr_4_1856) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_1856;
      ov := iv(0 downto 0);
      ptr_deref_1859_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1859_gather_scatter
    process(ptr_deref_1859_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1859_data_0;
      ov(15 downto 0) := iv;
      tmp21_1860 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1859_root_address_inst
    process(ptr_deref_1859_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1859_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1859_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_addr_0
    process(ptr_deref_1875_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1875_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1875_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_base_resize
    process(iNsTr_5_1872) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_1872;
      ov := iv(6 downto 0);
      ptr_deref_1875_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_gather_scatter
    process(ptr_deref_1875_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1875_data_0;
      ov(31 downto 0) := iv;
      tmp24_1876 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1875_root_address_inst
    process(ptr_deref_1875_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1875_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1875_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1892_addr_0
    process(ptr_deref_1892_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1892_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_1892_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1892_base_resize
    process(iNsTr_6_1889) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_1889;
      ov := iv(0 downto 0);
      ptr_deref_1892_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1892_gather_scatter
    process(ptr_deref_1892_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1892_data_0;
      ov(15 downto 0) := iv;
      tmp32_1893 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1892_root_address_inst
    process(ptr_deref_1892_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1892_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_1892_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1908_addr_0
    process(ptr_deref_1908_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1908_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1908_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1908_base_resize
    process(iNsTr_7_1905) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_1905;
      ov := iv(6 downto 0);
      ptr_deref_1908_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1908_gather_scatter
    process(ptr_deref_1908_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1908_data_0;
      ov(31 downto 0) := iv;
      tmp35_1909 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1908_root_address_inst
    process(ptr_deref_1908_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1908_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1908_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1920_addr_0
    process(ptr_deref_1920_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1920_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1920_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1920_base_resize
    process(iNsTr_8_1917) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_1917;
      ov := iv(6 downto 0);
      ptr_deref_1920_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1920_gather_scatter
    process(ptr_deref_1920_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1920_data_0;
      ov(31 downto 0) := iv;
      tmp44_1921 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1920_root_address_inst
    process(ptr_deref_1920_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1920_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1920_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1932_addr_0
    process(ptr_deref_1932_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1932_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1932_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1932_base_resize
    process(iNsTr_9_1929) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_1929;
      ov := iv(6 downto 0);
      ptr_deref_1932_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1932_gather_scatter
    process(ptr_deref_1932_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1932_data_0;
      ov(31 downto 0) := iv;
      tmp47_1933 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1932_root_address_inst
    process(ptr_deref_1932_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1932_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1932_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1944_addr_0
    process(ptr_deref_1944_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1944_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1944_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1944_base_resize
    process(iNsTr_10_1941) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_1941;
      ov := iv(6 downto 0);
      ptr_deref_1944_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1944_gather_scatter
    process(ptr_deref_1944_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1944_data_0;
      ov(31 downto 0) := iv;
      tmp87_1945 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1944_root_address_inst
    process(ptr_deref_1944_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1944_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1944_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2139_addr_0
    process(ptr_deref_2139_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2139_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2139_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2139_base_resize
    process(arrayidx_2136) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2136;
      ov := iv(13 downto 0);
      ptr_deref_2139_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2139_gather_scatter
    process(ptr_deref_2139_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2139_data_0;
      ov(63 downto 0) := iv;
      tmp57_2140 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2139_root_address_inst
    process(ptr_deref_2139_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2139_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2139_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_addr_0
    process(ptr_deref_2169_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_base_resize
    process(arrayidx62_2167) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx62_2167;
      ov := iv(13 downto 0);
      ptr_deref_2169_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_gather_scatter
    process(tmp57_2140) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp57_2140;
      ov(63 downto 0) := iv;
      ptr_deref_2169_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2169_root_address_inst
    process(ptr_deref_2169_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2169_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2169_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2188_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2187;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2188_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2188_branch_req_0,
          ack0 => if_stmt_2188_branch_ack_0,
          ack1 => if_stmt_2188_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2219_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp77_2218;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2219_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2219_branch_req_0,
          ack0 => if_stmt_2219_branch_ack_0,
          ack1 => if_stmt_2219_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2267_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp89_2266;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2267_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2267_branch_req_0,
          ack0 => if_stmt_2267_branch_ack_0,
          ack1 => if_stmt_2267_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2199_inst
    process(indvar_2082) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2082, type_cast_2198_wire_constant, tmp_var);
      indvarx_xnext_2200 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2207_inst
    process(input_dim1x_x1x_xph_1954) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_1954, type_cast_2206_wire_constant, tmp_var);
      inc_2208 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2230_inst
    process(input_dim0x_x2x_xph_1960) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_1960, type_cast_2229_wire_constant, tmp_var);
      inc81_2231 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1986_inst
    process(mul_1982, conv12_1972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_1982, conv12_1972, tmp_var);
      add_1987 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2001_inst
    process(mul23_1997, tmp24_1876) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul23_1997, tmp24_1876, tmp_var);
      add25_2002 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2016_inst
    process(mul34_2012, tmp35_1909) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul34_2012, tmp35_1909, tmp_var);
      add36_2017 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2033_inst
    process(sub40_2028) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub40_2028, type_cast_2032_wire_constant, tmp_var);
      sext_2034 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2054_inst
    process(sub28_2049) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub28_2049, type_cast_2053_wire_constant, tmp_var);
      sext103_2055 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2073_inst
    process(conv46_2043, mul50_2069) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv46_2043, mul50_2069, tmp_var);
      add51_2074 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2103_inst
    process(mul16_1992, conv9102_2099) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul16_1992, conv9102_2099, tmp_var);
      add17_2104 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2108_inst
    process(mul52_2079, conv9102_2099) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul52_2079, conv9102_2099, tmp_var);
      add53_2109 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2181_inst
    process(conv65_2176) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv65_2176, type_cast_2180_wire_constant, tmp_var);
      add66_2182 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2041_inst
    process(type_cast_2037_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2037_wire, type_cast_2040_wire_constant, tmp_var);
      ASHR_i32_i32_2041_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2062_inst
    process(type_cast_2058_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2058_wire, type_cast_2061_wire_constant, tmp_var);
      ASHR_i32_i32_2062_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2122_inst
    process(type_cast_2118_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2118_wire, type_cast_2121_wire_constant, tmp_var);
      ASHR_i32_i32_2122_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2153_inst
    process(type_cast_2149_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2149_wire, type_cast_2152_wire_constant, tmp_var);
      ASHR_i32_i32_2153_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2217_inst
    process(conv75_2213, tmp_1828) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv75_2213, tmp_1828, tmp_var);
      cmp77_2218 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2265_inst
    process(conv86_2261, div88_1951) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv86_2261, div88_1951, tmp_var);
      cmp89_2266 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1833_inst
    process(tmp_1828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1828, type_cast_1832_wire_constant, tmp_var);
      div_1834 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1950_inst
    process(tmp87_1945) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp87_1945, type_cast_1949_wire_constant, tmp_var);
      div88_1951 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2236_inst
    process(tmp_1828) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_1828, type_cast_2235_wire_constant, tmp_var);
      div83_2237 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2094_inst
    process(indvar_2082) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2082, type_cast_2093_wire_constant, tmp_var);
      input_dim2x_x1_2095 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1981_inst
    process(tmp_1828, conv15_1977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp_1828, conv15_1977, tmp_var);
      mul_1982 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1991_inst
    process(add_1987, tmp10_1850) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_1987, tmp10_1850, tmp_var);
      mul16_1992 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1996_inst
    process(conv22_1864, conv15_1977) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv22_1864, conv15_1977, tmp_var);
      mul23_1997 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2011_inst
    process(conv33_1897, conv12_1972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv33_1897, conv12_1972, tmp_var);
      mul34_2012 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2068_inst
    process(tmp47_1933, conv49_2064) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp47_1933, conv49_2064, tmp_var);
      mul50_2069 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2078_inst
    process(add51_2074, tmp44_1921) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add51_2074, tmp44_1921, tmp_var);
      mul52_2079 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2027_inst
    process(sub39_2022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub39_2022, type_cast_2026_wire_constant, tmp_var);
      sub40_2028 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2048_inst
    process(sub_2007) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2007, type_cast_2047_wire_constant, tmp_var);
      sub28_2049 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2114_inst
    process(add17_2104) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add17_2104, type_cast_2113_wire_constant, tmp_var);
      sext105_2115 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2145_inst
    process(add53_2109) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add53_2109, type_cast_2144_wire_constant, tmp_var);
      sext106_2146 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2006_inst
    process(add25_2002, conv27_1883) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add25_2002, conv27_1883, tmp_var);
      sub_2007 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2021_inst
    process(add36_2017, conv27_1883) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add36_2017, conv27_1883, tmp_var);
      sub39_2022 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2186_inst
    process(add66_2182, tmp10_1850) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add66_2182, tmp10_1850, tmp_var);
      cmp_2187 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_2134_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2133_scaled;
      array_obj_ref_2134_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2134_index_offset_req_0;
      array_obj_ref_2134_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2134_index_offset_req_1;
      array_obj_ref_2134_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_2165_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom61_2164_scaled;
      array_obj_ref_2165_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2165_index_offset_req_0;
      array_obj_ref_2165_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2165_index_offset_req_1;
      array_obj_ref_2165_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_1970_inst
    process(input_dim1x_x1x_xph_1954) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_1954, tmp_var);
      type_cast_1970_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1975_inst
    process(input_dim0x_x2x_xph_1960) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_1960, tmp_var);
      type_cast_1975_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2127_inst
    process(shr_2124) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2124, tmp_var);
      type_cast_2127_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2158_inst
    process(shr60_2155) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr60_2155, tmp_var);
      type_cast_2158_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2174_inst
    process(input_dim2x_x1_2095) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2095, tmp_var);
      type_cast_2174_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2211_inst
    process(inc_2208) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2208, tmp_var);
      type_cast_2211_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2259_inst
    process(input_dim0x_x0_2250) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_2250, tmp_var);
      type_cast_2259_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_1878_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_1878_load_0_req_0;
      LOAD_padding_1878_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_1878_load_0_req_1;
      LOAD_padding_1878_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_1878_word_address_0;
      LOAD_padding_1878_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1944_load_0 ptr_deref_1849_load_0 ptr_deref_1827_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1944_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1849_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1827_load_0_req_0;
      ptr_deref_1944_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1849_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1827_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1944_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1849_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1827_load_0_req_1;
      ptr_deref_1944_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1849_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1827_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1944_word_address_0 & ptr_deref_1849_word_address_0 & ptr_deref_1827_word_address_0;
      ptr_deref_1944_data_0 <= data_out(95 downto 64);
      ptr_deref_1849_data_0 <= data_out(63 downto 32);
      ptr_deref_1827_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1892_load_0 ptr_deref_1859_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1892_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1859_load_0_req_0;
      ptr_deref_1892_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1859_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1892_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1859_load_0_req_1;
      ptr_deref_1892_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1859_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1892_word_address_0 & ptr_deref_1859_word_address_0;
      ptr_deref_1892_data_0 <= data_out(31 downto 16);
      ptr_deref_1859_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1908_load_0 ptr_deref_1875_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1908_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1875_load_0_req_0;
      ptr_deref_1908_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1875_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1908_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1875_load_0_req_1;
      ptr_deref_1908_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1875_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1908_word_address_0 & ptr_deref_1875_word_address_0;
      ptr_deref_1908_data_0 <= data_out(63 downto 32);
      ptr_deref_1875_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_1920_load_0 ptr_deref_1932_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_1920_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1932_load_0_req_0;
      ptr_deref_1920_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1932_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_1920_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1932_load_0_req_1;
      ptr_deref_1920_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1932_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1920_word_address_0 & ptr_deref_1932_word_address_0;
      ptr_deref_1920_data_0 <= data_out(63 downto 32);
      ptr_deref_1932_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2139_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2139_load_0_req_0;
      ptr_deref_2139_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2139_load_0_req_1;
      ptr_deref_2139_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2139_word_address_0;
      ptr_deref_2139_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2169_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2169_store_0_req_0;
      ptr_deref_2169_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2169_store_0_req_1;
      ptr_deref_2169_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2169_word_address_0;
      data_in <= ptr_deref_2169_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block1_start_1814_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block1_start_1814_inst_req_0;
      RPIPE_Block1_start_1814_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block1_start_1814_inst_req_1;
      RPIPE_Block1_start_1814_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_1815 <= data_out(15 downto 0);
      Block1_start_read_0_gI: SplitGuardInterface generic map(name => "Block1_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block1_start_read_0: InputPortRevised -- 
        generic map ( name => "Block1_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block1_start_pipe_read_req(0),
          oack => Block1_start_pipe_read_ack(0),
          odata => Block1_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block1_done_2275_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block1_done_2275_inst_req_0;
      WPIPE_Block1_done_2275_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block1_done_2275_inst_req_1;
      WPIPE_Block1_done_2275_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_1815;
      Block1_done_write_0_gI: SplitGuardInterface generic map(name => "Block1_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block1_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block1_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block1_done_pipe_write_req(0),
          oack => Block1_done_pipe_write_ack(0),
          odata => Block1_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeB_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeC is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeC;
architecture convTransposeC_arch of convTransposeC is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeC_CP_6511_start: Boolean;
  signal convTransposeC_CP_6511_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal type_cast_2437_inst_req_0 : boolean;
  signal WPIPE_Block2_done_2724_inst_req_0 : boolean;
  signal type_cast_2431_inst_ack_1 : boolean;
  signal type_cast_2646_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2285_inst_ack_0 : boolean;
  signal RPIPE_Block2_start_2285_inst_ack_1 : boolean;
  signal type_cast_2646_inst_req_0 : boolean;
  signal ptr_deref_2298_load_0_req_1 : boolean;
  signal RPIPE_Block2_start_2285_inst_req_1 : boolean;
  signal WPIPE_Block2_done_2724_inst_ack_0 : boolean;
  signal type_cast_2437_inst_ack_0 : boolean;
  signal ptr_deref_2298_load_0_ack_1 : boolean;
  signal type_cast_2308_inst_req_1 : boolean;
  signal type_cast_2308_inst_req_0 : boolean;
  signal RPIPE_Block2_start_2285_inst_req_0 : boolean;
  signal type_cast_2308_inst_ack_0 : boolean;
  signal type_cast_2308_inst_ack_1 : boolean;
  signal ptr_deref_2298_load_0_ack_0 : boolean;
  signal phi_stmt_2425_req_1 : boolean;
  signal ptr_deref_2320_load_0_ack_0 : boolean;
  signal ptr_deref_2320_load_0_ack_1 : boolean;
  signal if_stmt_2659_branch_ack_1 : boolean;
  signal ptr_deref_2320_load_0_req_1 : boolean;
  signal if_stmt_2716_branch_ack_0 : boolean;
  signal ptr_deref_2320_load_0_req_0 : boolean;
  signal WPIPE_Block2_done_2724_inst_ack_1 : boolean;
  signal if_stmt_2716_branch_ack_1 : boolean;
  signal WPIPE_Block2_done_2724_inst_req_1 : boolean;
  signal ptr_deref_2332_load_0_req_0 : boolean;
  signal ptr_deref_2332_load_0_ack_0 : boolean;
  signal ptr_deref_2640_store_0_ack_1 : boolean;
  signal ptr_deref_2332_load_0_req_1 : boolean;
  signal ptr_deref_2332_load_0_ack_1 : boolean;
  signal phi_stmt_2432_ack_0 : boolean;
  signal phi_stmt_2432_req_0 : boolean;
  signal ptr_deref_2640_store_0_req_1 : boolean;
  signal type_cast_2431_inst_ack_0 : boolean;
  signal type_cast_2709_inst_ack_1 : boolean;
  signal type_cast_2709_inst_req_1 : boolean;
  signal type_cast_2431_inst_req_1 : boolean;
  signal type_cast_2709_inst_ack_0 : boolean;
  signal type_cast_2435_inst_ack_1 : boolean;
  signal type_cast_2709_inst_req_0 : boolean;
  signal type_cast_2435_inst_req_1 : boolean;
  signal ptr_deref_2298_load_0_req_0 : boolean;
  signal if_stmt_2659_branch_req_0 : boolean;
  signal ptr_deref_2342_load_0_req_0 : boolean;
  signal ptr_deref_2342_load_0_ack_0 : boolean;
  signal addr_of_2637_final_reg_ack_1 : boolean;
  signal if_stmt_2716_branch_req_0 : boolean;
  signal ptr_deref_2342_load_0_req_1 : boolean;
  signal ptr_deref_2342_load_0_ack_1 : boolean;
  signal phi_stmt_2425_ack_0 : boolean;
  signal type_cast_2692_inst_ack_1 : boolean;
  signal type_cast_2431_inst_req_0 : boolean;
  signal addr_of_2637_final_reg_req_1 : boolean;
  signal type_cast_2692_inst_req_1 : boolean;
  signal type_cast_2435_inst_ack_0 : boolean;
  signal type_cast_2346_inst_req_0 : boolean;
  signal type_cast_2435_inst_req_0 : boolean;
  signal type_cast_2346_inst_ack_0 : boolean;
  signal type_cast_2346_inst_req_1 : boolean;
  signal type_cast_2346_inst_ack_1 : boolean;
  signal ptr_deref_2640_store_0_ack_0 : boolean;
  signal ptr_deref_2358_load_0_req_0 : boolean;
  signal ptr_deref_2358_load_0_ack_0 : boolean;
  signal ptr_deref_2358_load_0_req_1 : boolean;
  signal ptr_deref_2358_load_0_ack_1 : boolean;
  signal ptr_deref_2640_store_0_req_0 : boolean;
  signal type_cast_2692_inst_ack_0 : boolean;
  signal type_cast_2692_inst_req_0 : boolean;
  signal LOAD_padding_2361_load_0_req_0 : boolean;
  signal LOAD_padding_2361_load_0_ack_0 : boolean;
  signal LOAD_padding_2361_load_0_req_1 : boolean;
  signal type_cast_2683_inst_ack_1 : boolean;
  signal LOAD_padding_2361_load_0_ack_1 : boolean;
  signal type_cast_2683_inst_req_1 : boolean;
  signal type_cast_2683_inst_ack_0 : boolean;
  signal type_cast_2683_inst_req_0 : boolean;
  signal phi_stmt_2432_req_1 : boolean;
  signal type_cast_2365_inst_req_0 : boolean;
  signal type_cast_2365_inst_ack_0 : boolean;
  signal addr_of_2637_final_reg_ack_0 : boolean;
  signal type_cast_2437_inst_ack_1 : boolean;
  signal type_cast_2365_inst_req_1 : boolean;
  signal phi_stmt_2425_req_0 : boolean;
  signal type_cast_2365_inst_ack_1 : boolean;
  signal addr_of_2637_final_reg_req_0 : boolean;
  signal type_cast_2646_inst_ack_1 : boolean;
  signal ptr_deref_2375_load_0_req_0 : boolean;
  signal ptr_deref_2375_load_0_ack_0 : boolean;
  signal type_cast_2646_inst_req_1 : boolean;
  signal ptr_deref_2375_load_0_req_1 : boolean;
  signal ptr_deref_2375_load_0_ack_1 : boolean;
  signal type_cast_2437_inst_req_1 : boolean;
  signal if_stmt_2659_branch_ack_0 : boolean;
  signal type_cast_2379_inst_req_0 : boolean;
  signal type_cast_2379_inst_ack_0 : boolean;
  signal type_cast_2379_inst_req_1 : boolean;
  signal type_cast_2379_inst_ack_1 : boolean;
  signal ptr_deref_2391_load_0_req_0 : boolean;
  signal ptr_deref_2391_load_0_ack_0 : boolean;
  signal ptr_deref_2391_load_0_req_1 : boolean;
  signal ptr_deref_2391_load_0_ack_1 : boolean;
  signal ptr_deref_2403_load_0_req_0 : boolean;
  signal ptr_deref_2403_load_0_ack_0 : boolean;
  signal ptr_deref_2403_load_0_req_1 : boolean;
  signal ptr_deref_2403_load_0_ack_1 : boolean;
  signal ptr_deref_2415_load_0_req_0 : boolean;
  signal ptr_deref_2415_load_0_ack_0 : boolean;
  signal ptr_deref_2415_load_0_req_1 : boolean;
  signal ptr_deref_2415_load_0_ack_1 : boolean;
  signal type_cast_2442_inst_req_0 : boolean;
  signal type_cast_2442_inst_ack_0 : boolean;
  signal type_cast_2442_inst_req_1 : boolean;
  signal type_cast_2442_inst_ack_1 : boolean;
  signal type_cast_2447_inst_req_0 : boolean;
  signal type_cast_2447_inst_ack_0 : boolean;
  signal type_cast_2447_inst_req_1 : boolean;
  signal type_cast_2447_inst_ack_1 : boolean;
  signal type_cast_2569_inst_req_0 : boolean;
  signal type_cast_2569_inst_ack_0 : boolean;
  signal type_cast_2569_inst_req_1 : boolean;
  signal type_cast_2569_inst_ack_1 : boolean;
  signal type_cast_2599_inst_req_0 : boolean;
  signal type_cast_2599_inst_ack_0 : boolean;
  signal type_cast_2599_inst_req_1 : boolean;
  signal type_cast_2599_inst_ack_1 : boolean;
  signal array_obj_ref_2605_index_offset_req_0 : boolean;
  signal array_obj_ref_2605_index_offset_ack_0 : boolean;
  signal array_obj_ref_2605_index_offset_req_1 : boolean;
  signal array_obj_ref_2605_index_offset_ack_1 : boolean;
  signal addr_of_2606_final_reg_req_0 : boolean;
  signal addr_of_2606_final_reg_ack_0 : boolean;
  signal addr_of_2606_final_reg_req_1 : boolean;
  signal addr_of_2606_final_reg_ack_1 : boolean;
  signal ptr_deref_2610_load_0_req_0 : boolean;
  signal ptr_deref_2610_load_0_ack_0 : boolean;
  signal ptr_deref_2610_load_0_req_1 : boolean;
  signal ptr_deref_2610_load_0_ack_1 : boolean;
  signal type_cast_2630_inst_req_0 : boolean;
  signal type_cast_2630_inst_ack_0 : boolean;
  signal type_cast_2630_inst_req_1 : boolean;
  signal type_cast_2630_inst_ack_1 : boolean;
  signal array_obj_ref_2636_index_offset_req_0 : boolean;
  signal array_obj_ref_2636_index_offset_ack_0 : boolean;
  signal array_obj_ref_2636_index_offset_req_1 : boolean;
  signal array_obj_ref_2636_index_offset_ack_1 : boolean;
  signal type_cast_2559_inst_req_0 : boolean;
  signal type_cast_2559_inst_ack_0 : boolean;
  signal type_cast_2559_inst_req_1 : boolean;
  signal type_cast_2559_inst_ack_1 : boolean;
  signal phi_stmt_2553_req_1 : boolean;
  signal phi_stmt_2553_req_0 : boolean;
  signal phi_stmt_2553_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeC_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeC_CP_6511_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeC_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeC_CP_6511_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeC_CP_6511: Block -- control-path 
    signal convTransposeC_CP_6511_elements: BooleanArray(92 downto 0);
    -- 
  begin -- 
    convTransposeC_CP_6511_elements(0) <= convTransposeC_CP_6511_start;
    convTransposeC_CP_6511_symbol <= convTransposeC_CP_6511_elements(70);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_2283/assign_stmt_2286/$entry
      -- CP-element group 0: 	 branch_block_stmt_2283/branch_block_stmt_2283__entry__
      -- CP-element group 0: 	 branch_block_stmt_2283/assign_stmt_2286__entry__
      -- CP-element group 0: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2283/$entry
      -- CP-element group 0: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Sample/rr
      -- 
    rr_6559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(0), ack => RPIPE_Block2_start_2285_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Update/cr
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_sample_completed_
      -- 
    ra_6560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2285_inst_ack_0, ack => convTransposeC_CP_6511_elements(1)); -- 
    cr_6564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(1), ack => RPIPE_Block2_start_2285_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	11 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	15 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	9 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	21 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	25 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2:  members (265) 
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2286__exit__
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2286/RPIPE_Block2_start_2285_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2286/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422__entry__
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/word_0/cr
      -- 
    ca_6565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block2_start_2285_inst_ack_1, ack => convTransposeC_CP_6511_elements(2)); -- 
    cr_6612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2298_load_0_req_1); -- 
    cr_6631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2308_inst_req_1); -- 
    cr_6676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2320_load_0_req_1); -- 
    rr_6665_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6665_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2320_load_0_req_0); -- 
    rr_6715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2332_load_0_req_0); -- 
    cr_6726_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6726_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2332_load_0_req_1); -- 
    rr_6601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2298_load_0_req_0); -- 
    rr_6765_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6765_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2342_load_0_req_0); -- 
    cr_6776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2342_load_0_req_1); -- 
    cr_6795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2346_inst_req_1); -- 
    rr_6829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2358_load_0_req_0); -- 
    cr_6840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2358_load_0_req_1); -- 
    rr_6862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => LOAD_padding_2361_load_0_req_0); -- 
    cr_6873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => LOAD_padding_2361_load_0_req_1); -- 
    cr_6892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2365_inst_req_1); -- 
    rr_6926_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6926_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2375_load_0_req_0); -- 
    cr_6937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2375_load_0_req_1); -- 
    cr_6956_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_6956_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => type_cast_2379_inst_req_1); -- 
    rr_6990_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6990_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2391_load_0_req_0); -- 
    cr_7001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2391_load_0_req_1); -- 
    rr_7040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2403_load_0_req_0); -- 
    cr_7051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2403_load_0_req_1); -- 
    rr_7090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2415_load_0_req_0); -- 
    cr_7101_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7101_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(2), ack => ptr_deref_2415_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Sample/word_access_start/word_0/ra
      -- 
    ra_6602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2298_load_0_ack_0, ack => convTransposeC_CP_6511_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/ptr_deref_2298_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/ptr_deref_2298_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/ptr_deref_2298_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2298_Update/ptr_deref_2298_Merge/$entry
      -- 
    ca_6613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2298_load_0_ack_1, ack => convTransposeC_CP_6511_elements(4)); -- 
    rr_6626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(4), ack => type_cast_2308_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Sample/ra
      -- 
    ra_6627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_0, ack => convTransposeC_CP_6511_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2308_Update/ca
      -- 
    ca_6632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2308_inst_ack_1, ack => convTransposeC_CP_6511_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/word_0/ra
      -- CP-element group 7: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Sample/$exit
      -- 
    ra_6666_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2320_load_0_ack_0, ack => convTransposeC_CP_6511_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	31 
    -- CP-element group 8:  members (9) 
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/ptr_deref_2320_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/ptr_deref_2320_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/ptr_deref_2320_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/ptr_deref_2320_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2320_Update/$exit
      -- 
    ca_6677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2320_load_0_ack_1, ack => convTransposeC_CP_6511_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	2 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/word_0/$exit
      -- CP-element group 9: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/word_0/ra
      -- CP-element group 9: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Sample/word_access_start/$exit
      -- 
    ra_6716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2332_load_0_ack_0, ack => convTransposeC_CP_6511_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	31 
    -- CP-element group 10:  members (9) 
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/$exit
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/word_0/$exit
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/word_access_complete/word_0/ca
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/ptr_deref_2332_Merge/$entry
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/ptr_deref_2332_Merge/$exit
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/ptr_deref_2332_Merge/merge_req
      -- CP-element group 10: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2332_Update/ptr_deref_2332_Merge/merge_ack
      -- 
    ca_6727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2332_load_0_ack_1, ack => convTransposeC_CP_6511_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Sample/word_access_start/word_0/ra
      -- 
    ra_6766_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2342_load_0_ack_0, ack => convTransposeC_CP_6511_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (12) 
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/ptr_deref_2342_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/ptr_deref_2342_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/ptr_deref_2342_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2342_Update/ptr_deref_2342_Merge/merge_ack
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Sample/rr
      -- 
    ca_6777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2342_load_0_ack_1, ack => convTransposeC_CP_6511_elements(12)); -- 
    rr_6790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(12), ack => type_cast_2346_inst_req_0); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Sample/ra
      -- 
    ra_6791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_0, ack => convTransposeC_CP_6511_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	31 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2346_Update/ca
      -- 
    ca_6796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2346_inst_ack_1, ack => convTransposeC_CP_6511_elements(14)); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (5) 
      -- CP-element group 15: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/$exit
      -- CP-element group 15: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/word_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Sample/word_access_start/word_0/ra
      -- 
    ra_6830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_load_0_ack_0, ack => convTransposeC_CP_6511_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (9) 
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/$exit
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/word_access_complete/word_0/ca
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/ptr_deref_2358_Merge/$entry
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/ptr_deref_2358_Merge/$exit
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/ptr_deref_2358_Merge/merge_req
      -- CP-element group 16: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2358_Update/ptr_deref_2358_Merge/merge_ack
      -- 
    ca_6841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2358_load_0_ack_1, ack => convTransposeC_CP_6511_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Sample/word_access_start/word_0/ra
      -- 
    ra_6863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2361_load_0_ack_0, ack => convTransposeC_CP_6511_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (12) 
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/LOAD_padding_2361_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/LOAD_padding_2361_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/LOAD_padding_2361_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/LOAD_padding_2361_Update/LOAD_padding_2361_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Sample/rr
      -- 
    ca_6874_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2361_load_0_ack_1, ack => convTransposeC_CP_6511_elements(18)); -- 
    rr_6887_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6887_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(18), ack => type_cast_2365_inst_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Sample/ra
      -- 
    ra_6888_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_0, ack => convTransposeC_CP_6511_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	31 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2365_Update/ca
      -- 
    ca_6893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2365_inst_ack_1, ack => convTransposeC_CP_6511_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	2 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Sample/word_access_start/word_0/ra
      -- 
    ra_6927_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2375_load_0_ack_0, ack => convTransposeC_CP_6511_elements(21)); -- 
    -- CP-element group 22:  transition  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (12) 
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/word_access_complete/word_0/ca
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/ptr_deref_2375_Merge/$entry
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/ptr_deref_2375_Merge/$exit
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/ptr_deref_2375_Merge/merge_req
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2375_Update/ptr_deref_2375_Merge/merge_ack
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Sample/rr
      -- 
    ca_6938_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2375_load_0_ack_1, ack => convTransposeC_CP_6511_elements(22)); -- 
    rr_6951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_6951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(22), ack => type_cast_2379_inst_req_0); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Sample/ra
      -- 
    ra_6952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2379_inst_ack_0, ack => convTransposeC_CP_6511_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	31 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/type_cast_2379_Update/ca
      -- 
    ca_6957_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2379_inst_ack_1, ack => convTransposeC_CP_6511_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	2 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (5) 
      -- CP-element group 25: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/$exit
      -- CP-element group 25: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Sample/word_access_start/word_0/ra
      -- 
    ra_6991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2391_load_0_ack_0, ack => convTransposeC_CP_6511_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	31 
    -- CP-element group 26:  members (9) 
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/$exit
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/word_0/$exit
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/word_access_complete/word_0/ca
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/ptr_deref_2391_Merge/$entry
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/ptr_deref_2391_Merge/$exit
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/ptr_deref_2391_Merge/merge_req
      -- CP-element group 26: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2391_Update/ptr_deref_2391_Merge/merge_ack
      -- 
    ca_7002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2391_load_0_ack_1, ack => convTransposeC_CP_6511_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Sample/word_access_start/word_0/ra
      -- 
    ra_7041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2403_load_0_ack_0, ack => convTransposeC_CP_6511_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	31 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/ptr_deref_2403_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/ptr_deref_2403_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/ptr_deref_2403_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2403_Update/ptr_deref_2403_Merge/merge_ack
      -- 
    ca_7052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2403_load_0_ack_1, ack => convTransposeC_CP_6511_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Sample/word_access_start/word_0/ra
      -- 
    ra_7091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2415_load_0_ack_0, ack => convTransposeC_CP_6511_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	31 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/ptr_deref_2415_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/ptr_deref_2415_Merge/$exit
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/ptr_deref_2415_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/ptr_deref_2415_Update/ptr_deref_2415_Merge/merge_ack
      -- 
    ca_7102_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2415_load_0_ack_1, ack => convTransposeC_CP_6511_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	30 
    -- CP-element group 31: 	14 
    -- CP-element group 31: 	8 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	20 
    -- CP-element group 31: 	10 
    -- CP-element group 31: 	24 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	28 
    -- CP-element group 31: 	6 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	71 
    -- CP-element group 31: 	72 
    -- CP-element group 31: 	73 
    -- CP-element group 31:  members (14) 
      -- CP-element group 31: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422__exit__
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter
      -- CP-element group 31: 	 branch_block_stmt_2283/assign_stmt_2295_to_assign_stmt_2422/$exit
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Update/cr
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Sample/rr
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/$entry
      -- CP-element group 31: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$entry
      -- 
    cr_7524_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7524_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(31), ack => type_cast_2435_inst_req_1); -- 
    rr_7519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(31), ack => type_cast_2435_inst_req_0); -- 
    convTransposeC_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(30) & convTransposeC_CP_6511_elements(14) & convTransposeC_CP_6511_elements(8) & convTransposeC_CP_6511_elements(16) & convTransposeC_CP_6511_elements(20) & convTransposeC_CP_6511_elements(10) & convTransposeC_CP_6511_elements(24) & convTransposeC_CP_6511_elements(26) & convTransposeC_CP_6511_elements(28) & convTransposeC_CP_6511_elements(6);
      gj_convTransposeC_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	86 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Sample/ra
      -- 
    ra_7119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_0, ack => convTransposeC_CP_6511_elements(32)); -- 
    -- CP-element group 33:  transition  input  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	86 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	36 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Update/ca
      -- 
    ca_7124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2442_inst_ack_1, ack => convTransposeC_CP_6511_elements(33)); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	86 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Sample/ra
      -- 
    ra_7133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_0, ack => convTransposeC_CP_6511_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	86 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Update/ca
      -- 
    ca_7138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2447_inst_ack_1, ack => convTransposeC_CP_6511_elements(35)); -- 
    -- CP-element group 36:  join  transition  place  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	33 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	90 
    -- CP-element group 36:  members (6) 
      -- CP-element group 36: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550__exit__
      -- CP-element group 36: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 36: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/$exit
      -- CP-element group 36: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/$entry
      -- CP-element group 36: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$entry
      -- 
    convTransposeC_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(35) & convTransposeC_CP_6511_elements(33);
      gj_convTransposeC_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Sample/ra
      -- 
    ra_7150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2569_inst_ack_0, ack => convTransposeC_CP_6511_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  output  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	92 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	47 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (9) 
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Update/ca
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Sample/rr
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Sample/rr
      -- 
    ca_7155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2569_inst_ack_1, ack => convTransposeC_CP_6511_elements(38)); -- 
    rr_7163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(38), ack => type_cast_2599_inst_req_0); -- 
    rr_7273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(38), ack => type_cast_2630_inst_req_0); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Sample/ra
      -- 
    ra_7164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_0, ack => convTransposeC_CP_6511_elements(39)); -- 
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	92 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (16) 
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_resized_1
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_scaled_1
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_computed_1
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_resize_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_resize_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_resize_1/index_resize_req
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_resize_1/index_resize_ack
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_scale_1/$entry
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_scale_1/$exit
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_scale_1/scale_rename_req
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_index_scale_1/scale_rename_ack
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Sample/req
      -- 
    ca_7169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2599_inst_ack_1, ack => convTransposeC_CP_6511_elements(40)); -- 
    req_7194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(40), ack => array_obj_ref_2605_index_offset_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_sample_complete
      -- CP-element group 41: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Sample/ack
      -- 
    ack_7195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2605_index_offset_ack_0, ack => convTransposeC_CP_6511_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	92 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (11) 
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_root_address_calculated
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_offset_calculated
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Update/ack
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_base_plus_offset/$entry
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_base_plus_offset/$exit
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_base_plus_offset/sum_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_base_plus_offset/sum_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_request/$entry
      -- CP-element group 42: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_request/req
      -- 
    ack_7200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2605_index_offset_ack_1, ack => convTransposeC_CP_6511_elements(42)); -- 
    req_7209_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7209_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(42), ack => addr_of_2606_final_reg_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_request/$exit
      -- CP-element group 43: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_request/ack
      -- 
    ack_7210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2606_final_reg_ack_0, ack => convTransposeC_CP_6511_elements(43)); -- 
    -- CP-element group 44:  join  fork  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	92 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (24) 
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_complete/$exit
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_complete/ack
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_word_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_address_resized
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_addr_resize/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_addr_resize/$exit
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_addr_resize/base_resize_req
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_addr_resize/base_resize_ack
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_word_addrgen/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_word_addrgen/$exit
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_word_addrgen/root_register_req
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_word_addrgen/root_register_ack
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/word_0/$entry
      -- CP-element group 44: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/word_0/rr
      -- 
    ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2606_final_reg_ack_1, ack => convTransposeC_CP_6511_elements(44)); -- 
    rr_7248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(44), ack => ptr_deref_2610_load_0_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (5) 
      -- CP-element group 45: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/$exit
      -- CP-element group 45: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/$exit
      -- CP-element group 45: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/word_0/$exit
      -- CP-element group 45: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Sample/word_access_start/word_0/ra
      -- 
    ra_7249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2610_load_0_ack_0, ack => convTransposeC_CP_6511_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	92 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	53 
    -- CP-element group 46:  members (9) 
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/$exit
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/word_0/$exit
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/word_0/ca
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/ptr_deref_2610_Merge/$entry
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/ptr_deref_2610_Merge/$exit
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/ptr_deref_2610_Merge/merge_req
      -- CP-element group 46: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/ptr_deref_2610_Merge/merge_ack
      -- 
    ca_7260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2610_load_0_ack_1, ack => convTransposeC_CP_6511_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	38 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Sample/ra
      -- 
    ra_7274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_0, ack => convTransposeC_CP_6511_elements(47)); -- 
    -- CP-element group 48:  transition  input  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	92 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (16) 
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Update/ca
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_resized_1
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_scaled_1
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_computed_1
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_resize_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_resize_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_resize_1/index_resize_req
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_resize_1/index_resize_ack
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_scale_1/$entry
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_scale_1/$exit
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_scale_1/scale_rename_req
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_index_scale_1/scale_rename_ack
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Sample/req
      -- 
    ca_7279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2630_inst_ack_1, ack => convTransposeC_CP_6511_elements(48)); -- 
    req_7304_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7304_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(48), ack => array_obj_ref_2636_index_offset_req_0); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_sample_complete
      -- CP-element group 49: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Sample/ack
      -- 
    ack_7305_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2636_index_offset_ack_0, ack => convTransposeC_CP_6511_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	92 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (11) 
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_request/req
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_request/$entry
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_root_address_calculated
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_offset_calculated
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Update/ack
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/$entry
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/$exit
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/sum_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_base_plus_offset/sum_rename_ack
      -- 
    ack_7310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2636_index_offset_ack_1, ack => convTransposeC_CP_6511_elements(50)); -- 
    req_7319_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7319_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(50), ack => addr_of_2637_final_reg_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_request/ack
      -- CP-element group 51: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_request/$exit
      -- CP-element group 51: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_sample_completed_
      -- 
    ack_7320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2637_final_reg_ack_0, ack => convTransposeC_CP_6511_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	92 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (19) 
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_word_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_complete/ack
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_complete/$exit
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_word_addrgen/root_register_ack
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_word_addrgen/root_register_req
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_word_addrgen/$exit
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_word_addrgen/$entry
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_addr_resize/base_resize_ack
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_addr_resize/base_resize_req
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_addr_resize/$exit
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_addr_resize/$entry
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_base_address_resized
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_update_completed_
      -- 
    ack_7325_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2637_final_reg_ack_1, ack => convTransposeC_CP_6511_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: 	46 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/ptr_deref_2640_Split/$exit
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/ptr_deref_2640_Split/$entry
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/word_0/rr
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/word_0/$entry
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/$entry
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/ptr_deref_2640_Split/split_ack
      -- CP-element group 53: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/ptr_deref_2640_Split/split_req
      -- 
    rr_7363_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7363_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(53), ack => ptr_deref_2640_store_0_req_0); -- 
    convTransposeC_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(52) & convTransposeC_CP_6511_elements(46);
      gj_convTransposeC_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (5) 
      -- CP-element group 54: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/word_0/ra
      -- CP-element group 54: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/word_0/$exit
      -- CP-element group 54: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Sample/word_access_start/$exit
      -- 
    ra_7364_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_store_0_ack_0, ack => convTransposeC_CP_6511_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	92 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	58 
    -- CP-element group 55:  members (5) 
      -- CP-element group 55: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/word_0/ca
      -- CP-element group 55: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/word_0/$exit
      -- CP-element group 55: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/$exit
      -- CP-element group 55: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/$exit
      -- 
    ca_7375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2640_store_0_ack_1, ack => convTransposeC_CP_6511_elements(55)); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	92 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_sample_completed_
      -- 
    ra_7384_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2646_inst_ack_0, ack => convTransposeC_CP_6511_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	92 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Update/ca
      -- 
    ca_7389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2646_inst_ack_1, ack => convTransposeC_CP_6511_elements(57)); -- 
    -- CP-element group 58:  branch  join  transition  place  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	41 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	55 
    -- CP-element group 58: 	49 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (10) 
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659__entry__
      -- CP-element group 58: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658__exit__
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_else_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2283/R_cmp_2660_place
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_if_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_eval_test/branch_req
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_eval_test/$exit
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_eval_test/$entry
      -- CP-element group 58: 	 branch_block_stmt_2283/if_stmt_2659_dead_link/$entry
      -- CP-element group 58: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/$exit
      -- 
    branch_req_7397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(58), ack => if_stmt_2659_branch_req_0); -- 
    convTransposeC_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(41) & convTransposeC_CP_6511_elements(57) & convTransposeC_CP_6511_elements(55) & convTransposeC_CP_6511_elements(49);
      gj_convTransposeC_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	87 
    -- CP-element group 59: 	88 
    -- CP-element group 59:  members (24) 
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody
      -- CP-element group 59: 	 branch_block_stmt_2283/assign_stmt_2671__exit__
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/merge_stmt_2665__exit__
      -- CP-element group 59: 	 branch_block_stmt_2283/assign_stmt_2671__entry__
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/if_stmt_2659_if_link/if_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_2283/whilex_xbody_ifx_xthen
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/if_stmt_2659_if_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/assign_stmt_2671/$exit
      -- CP-element group 59: 	 branch_block_stmt_2283/assign_stmt_2671/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Update/cr
      -- CP-element group 59: 	 branch_block_stmt_2283/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 59: 	 branch_block_stmt_2283/merge_stmt_2665_PhiReqMerge
      -- CP-element group 59: 	 branch_block_stmt_2283/merge_stmt_2665_PhiAck/$entry
      -- CP-element group 59: 	 branch_block_stmt_2283/merge_stmt_2665_PhiAck/$exit
      -- CP-element group 59: 	 branch_block_stmt_2283/merge_stmt_2665_PhiAck/dummy
      -- 
    if_choice_transition_7402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2659_branch_ack_1, ack => convTransposeC_CP_6511_elements(59)); -- 
    rr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7600_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(59), ack => type_cast_2559_inst_req_0); -- 
    cr_7605_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7605_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(59), ack => type_cast_2559_inst_req_1); -- 
    -- CP-element group 60:  fork  transition  place  input  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60: 	64 
    -- CP-element group 60: 	66 
    -- CP-element group 60:  members (24) 
      -- CP-element group 60: 	 branch_block_stmt_2283/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715__entry__
      -- CP-element group 60: 	 branch_block_stmt_2283/merge_stmt_2673__exit__
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2283/whilex_xbody_ifx_xelse
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Update/cr
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Sample/rr
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Sample/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_update_start_
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/if_stmt_2659_else_link/else_choice_transition
      -- CP-element group 60: 	 branch_block_stmt_2283/if_stmt_2659_else_link/$exit
      -- CP-element group 60: 	 branch_block_stmt_2283/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_2283/merge_stmt_2673_PhiReqMerge
      -- CP-element group 60: 	 branch_block_stmt_2283/merge_stmt_2673_PhiAck/$entry
      -- CP-element group 60: 	 branch_block_stmt_2283/merge_stmt_2673_PhiAck/$exit
      -- CP-element group 60: 	 branch_block_stmt_2283/merge_stmt_2673_PhiAck/dummy
      -- 
    else_choice_transition_7406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2659_branch_ack_0, ack => convTransposeC_CP_6511_elements(60)); -- 
    cr_7455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2709_inst_req_1); -- 
    cr_7441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2692_inst_req_1); -- 
    cr_7427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2683_inst_req_1); -- 
    rr_7422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(60), ack => type_cast_2683_inst_req_0); -- 
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Sample/ra
      -- CP-element group 61: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_sample_completed_
      -- 
    ra_7423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2683_inst_ack_0, ack => convTransposeC_CP_6511_elements(61)); -- 
    -- CP-element group 62:  transition  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (6) 
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Update/ca
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2683_update_completed_
      -- 
    ca_7428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2683_inst_ack_1, ack => convTransposeC_CP_6511_elements(62)); -- 
    rr_7436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(62), ack => type_cast_2692_inst_req_0); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Sample/ra
      -- CP-element group 63: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_sample_completed_
      -- 
    ra_7437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_0, ack => convTransposeC_CP_6511_elements(63)); -- 
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Sample/rr
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2692_update_completed_
      -- 
    ca_7442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2692_inst_ack_1, ack => convTransposeC_CP_6511_elements(64)); -- 
    rr_7450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(64), ack => type_cast_2709_inst_req_0); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Sample/ra
      -- CP-element group 65: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Sample/$exit
      -- CP-element group 65: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_sample_completed_
      -- 
    ra_7451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_0, ack => convTransposeC_CP_6511_elements(65)); -- 
    -- CP-element group 66:  branch  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	60 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (13) 
      -- CP-element group 66: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715__exit__
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716__entry__
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_else_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2283/R_cmp87_2717_place
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_eval_test/$exit
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_eval_test/$entry
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_dead_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Update/ca
      -- CP-element group 66: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_Update/$exit
      -- CP-element group 66: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/type_cast_2709_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_if_link/$entry
      -- CP-element group 66: 	 branch_block_stmt_2283/if_stmt_2716_eval_test/branch_req
      -- CP-element group 66: 	 branch_block_stmt_2283/assign_stmt_2679_to_assign_stmt_2715/$exit
      -- 
    ca_7456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2709_inst_ack_1, ack => convTransposeC_CP_6511_elements(66)); -- 
    branch_req_7464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_7464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(66), ack => if_stmt_2716_branch_req_0); -- 
    -- CP-element group 67:  merge  transition  place  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (15) 
      -- CP-element group 67: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Sample/req
      -- CP-element group 67: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_2283/merge_stmt_2722__exit__
      -- CP-element group 67: 	 branch_block_stmt_2283/assign_stmt_2726__entry__
      -- CP-element group 67: 	 branch_block_stmt_2283/ifx_xelse_whilex_xend
      -- CP-element group 67: 	 branch_block_stmt_2283/assign_stmt_2726/$entry
      -- CP-element group 67: 	 branch_block_stmt_2283/if_stmt_2716_if_link/if_choice_transition
      -- CP-element group 67: 	 branch_block_stmt_2283/if_stmt_2716_if_link/$exit
      -- CP-element group 67: 	 branch_block_stmt_2283/ifx_xelse_whilex_xend_PhiReq/$entry
      -- CP-element group 67: 	 branch_block_stmt_2283/ifx_xelse_whilex_xend_PhiReq/$exit
      -- CP-element group 67: 	 branch_block_stmt_2283/merge_stmt_2722_PhiReqMerge
      -- CP-element group 67: 	 branch_block_stmt_2283/merge_stmt_2722_PhiAck/$entry
      -- CP-element group 67: 	 branch_block_stmt_2283/merge_stmt_2722_PhiAck/$exit
      -- CP-element group 67: 	 branch_block_stmt_2283/merge_stmt_2722_PhiAck/dummy
      -- 
    if_choice_transition_7469_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2716_branch_ack_1, ack => convTransposeC_CP_6511_elements(67)); -- 
    req_7486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(67), ack => WPIPE_Block2_done_2724_inst_req_0); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	76 
    -- CP-element group 68: 	77 
    -- CP-element group 68: 	79 
    -- CP-element group 68: 	80 
    -- CP-element group 68:  members (20) 
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/if_stmt_2716_else_link/$exit
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/if_stmt_2716_else_link/else_choice_transition
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/$entry
      -- 
    else_choice_transition_7473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2716_branch_ack_0, ack => convTransposeC_CP_6511_elements(68)); -- 
    rr_7568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2437_inst_req_0); -- 
    cr_7550_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7550_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2431_inst_req_1); -- 
    rr_7545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2431_inst_req_0); -- 
    cr_7573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(68), ack => type_cast_2437_inst_req_1); -- 
    -- CP-element group 69:  transition  input  output  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (6) 
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Sample/ack
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_update_start_
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Update/req
      -- 
    ack_7487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2724_inst_ack_0, ack => convTransposeC_CP_6511_elements(69)); -- 
    req_7491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(69), ack => WPIPE_Block2_done_2724_inst_req_1); -- 
    -- CP-element group 70:  transition  place  input  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (16) 
      -- CP-element group 70: 	 branch_block_stmt_2283/$exit
      -- CP-element group 70: 	 $exit
      -- CP-element group 70: 	 branch_block_stmt_2283/branch_block_stmt_2283__exit__
      -- CP-element group 70: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2283/assign_stmt_2726/$exit
      -- CP-element group 70: 	 branch_block_stmt_2283/assign_stmt_2726__exit__
      -- CP-element group 70: 	 branch_block_stmt_2283/return__
      -- CP-element group 70: 	 branch_block_stmt_2283/merge_stmt_2728__exit__
      -- CP-element group 70: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Update/ack
      -- CP-element group 70: 	 branch_block_stmt_2283/assign_stmt_2726/WPIPE_Block2_done_2724_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2283/return___PhiReq/$entry
      -- CP-element group 70: 	 branch_block_stmt_2283/return___PhiReq/$exit
      -- CP-element group 70: 	 branch_block_stmt_2283/merge_stmt_2728_PhiReqMerge
      -- CP-element group 70: 	 branch_block_stmt_2283/merge_stmt_2728_PhiAck/$entry
      -- CP-element group 70: 	 branch_block_stmt_2283/merge_stmt_2728_PhiAck/$exit
      -- CP-element group 70: 	 branch_block_stmt_2283/merge_stmt_2728_PhiAck/dummy
      -- 
    ack_7492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block2_done_2724_inst_ack_1, ack => convTransposeC_CP_6511_elements(70)); -- 
    -- CP-element group 71:  transition  output  delay-element  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	31 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	75 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_req
      -- CP-element group 71: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2429_konst_delay_trans
      -- CP-element group 71: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$exit
      -- CP-element group 71: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/$exit
      -- 
    phi_stmt_2425_req_7503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2425_req_7503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(71), ack => phi_stmt_2425_req_0); -- 
    -- Element group convTransposeC_CP_6511_elements(71) is a control-delay.
    cp_element_71_delay: control_delay_element  generic map(name => " 71_delay", delay_value => 1)  port map(req => convTransposeC_CP_6511_elements(31), ack => convTransposeC_CP_6511_elements(71), clk => clk, reset =>reset);
    -- CP-element group 72:  transition  input  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	31 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (2) 
      -- CP-element group 72: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Sample/$exit
      -- 
    ra_7520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2435_inst_ack_0, ack => convTransposeC_CP_6511_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	31 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (2) 
      -- CP-element group 73: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Update/ca
      -- CP-element group 73: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/Update/$exit
      -- 
    ca_7525_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2435_inst_ack_1, ack => convTransposeC_CP_6511_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	75 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_req
      -- CP-element group 74: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/SplitProtocol/$exit
      -- CP-element group 74: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2435/$exit
      -- CP-element group 74: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/$exit
      -- CP-element group 74: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/$exit
      -- 
    phi_stmt_2432_req_7526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2432_req_7526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(74), ack => phi_stmt_2432_req_0); -- 
    convTransposeC_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(72) & convTransposeC_CP_6511_elements(73);
      gj_convTransposeC_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	71 
    -- CP-element group 75: 	74 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	83 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2283/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(71) & convTransposeC_CP_6511_elements(74);
      gj_convTransposeC_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	68 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Sample/$exit
      -- 
    ra_7546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_0, ack => convTransposeC_CP_6511_elements(76)); -- 
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	68 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/ca
      -- CP-element group 77: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/Update/$exit
      -- 
    ca_7551_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2431_inst_ack_1, ack => convTransposeC_CP_6511_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	82 
    -- CP-element group 78:  members (5) 
      -- CP-element group 78: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/$exit
      -- CP-element group 78: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_req
      -- CP-element group 78: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/$exit
      -- CP-element group 78: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/SplitProtocol/$exit
      -- CP-element group 78: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2425/phi_stmt_2425_sources/type_cast_2431/$exit
      -- 
    phi_stmt_2425_req_7552_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2425_req_7552_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(78), ack => phi_stmt_2425_req_1); -- 
    convTransposeC_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(76) & convTransposeC_CP_6511_elements(77);
      gj_convTransposeC_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	68 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Sample/$exit
      -- 
    ra_7569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_0, ack => convTransposeC_CP_6511_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	68 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Update/ca
      -- CP-element group 80: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/Update/$exit
      -- 
    ca_7574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2437_inst_ack_1, ack => convTransposeC_CP_6511_elements(80)); -- 
    -- CP-element group 81:  join  transition  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/$exit
      -- CP-element group 81: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/SplitProtocol/$exit
      -- CP-element group 81: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/type_cast_2437/$exit
      -- CP-element group 81: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_req
      -- CP-element group 81: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/phi_stmt_2432/phi_stmt_2432_sources/$exit
      -- 
    phi_stmt_2432_req_7575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2432_req_7575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(81), ack => phi_stmt_2432_req_1); -- 
    convTransposeC_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(79) & convTransposeC_CP_6511_elements(80);
      gj_convTransposeC_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  join  transition  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	78 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	83 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_2283/ifx_xelse_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeC_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(78) & convTransposeC_CP_6511_elements(81);
      gj_convTransposeC_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  merge  fork  transition  place  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	75 
    -- CP-element group 83: 	82 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2283/merge_stmt_2424_PhiAck/$entry
      -- CP-element group 83: 	 branch_block_stmt_2283/merge_stmt_2424_PhiReqMerge
      -- 
    convTransposeC_CP_6511_elements(83) <= OrReduce(convTransposeC_CP_6511_elements(75) & convTransposeC_CP_6511_elements(82));
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (1) 
      -- CP-element group 84: 	 branch_block_stmt_2283/merge_stmt_2424_PhiAck/phi_stmt_2425_ack
      -- 
    phi_stmt_2425_ack_7580_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2425_ack_0, ack => convTransposeC_CP_6511_elements(84)); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	86 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_2283/merge_stmt_2424_PhiAck/phi_stmt_2432_ack
      -- 
    phi_stmt_2432_ack_7581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2432_ack_0, ack => convTransposeC_CP_6511_elements(85)); -- 
    -- CP-element group 86:  join  fork  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: 	85 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	34 
    -- CP-element group 86: 	35 
    -- CP-element group 86: 	32 
    -- CP-element group 86: 	33 
    -- CP-element group 86:  members (16) 
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550__entry__
      -- CP-element group 86: 	 branch_block_stmt_2283/merge_stmt_2424__exit__
      -- CP-element group 86: 	 branch_block_stmt_2283/merge_stmt_2424_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/$entry
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2442_Update/cr
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_sample_start_
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_update_start_
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_2283/assign_stmt_2443_to_assign_stmt_2550/type_cast_2447_Update/cr
      -- 
    rr_7118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2442_inst_req_0); -- 
    cr_7123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2442_inst_req_1); -- 
    rr_7132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2447_inst_req_0); -- 
    cr_7137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(86), ack => type_cast_2447_inst_req_1); -- 
    convTransposeC_cp_element_group_86: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_86"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(84) & convTransposeC_CP_6511_elements(85);
      gj_convTransposeC_cp_element_group_86 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(86), clk => clk, reset => reset); --
    end block;
    -- CP-element group 87:  transition  input  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	59 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (2) 
      -- CP-element group 87: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Sample/$exit
      -- CP-element group 87: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Sample/ra
      -- 
    ra_7601_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_0, ack => convTransposeC_CP_6511_elements(87)); -- 
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	59 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Update/$exit
      -- CP-element group 88: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/Update/ca
      -- 
    ca_7606_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2559_inst_ack_1, ack => convTransposeC_CP_6511_elements(88)); -- 
    -- CP-element group 89:  join  transition  output  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (6) 
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$exit
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/$exit
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/$exit
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2559/SplitProtocol/$exit
      -- CP-element group 89: 	 branch_block_stmt_2283/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_req
      -- 
    phi_stmt_2553_req_7607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2553_req_7607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(89), ack => phi_stmt_2553_req_1); -- 
    convTransposeC_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeC_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeC_CP_6511_elements(87) & convTransposeC_CP_6511_elements(88);
      gj_convTransposeC_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeC_CP_6511_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  transition  output  delay-element  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	36 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (5) 
      -- CP-element group 90: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 90: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/$exit
      -- CP-element group 90: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/$exit
      -- CP-element group 90: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_sources/type_cast_2557_konst_delay_trans
      -- CP-element group 90: 	 branch_block_stmt_2283/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_2553/phi_stmt_2553_req
      -- 
    phi_stmt_2553_req_7618_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2553_req_7618_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(90), ack => phi_stmt_2553_req_0); -- 
    -- Element group convTransposeC_CP_6511_elements(90) is a control-delay.
    cp_element_90_delay: control_delay_element  generic map(name => " 90_delay", delay_value => 1)  port map(req => convTransposeC_CP_6511_elements(36), ack => convTransposeC_CP_6511_elements(90), clk => clk, reset =>reset);
    -- CP-element group 91:  merge  transition  place  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (2) 
      -- CP-element group 91: 	 branch_block_stmt_2283/merge_stmt_2552_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_2283/merge_stmt_2552_PhiAck/$entry
      -- 
    convTransposeC_CP_6511_elements(91) <= OrReduce(convTransposeC_CP_6511_elements(89) & convTransposeC_CP_6511_elements(90));
    -- CP-element group 92:  fork  transition  place  input  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	44 
    -- CP-element group 92: 	42 
    -- CP-element group 92: 	48 
    -- CP-element group 92: 	37 
    -- CP-element group 92: 	38 
    -- CP-element group 92: 	40 
    -- CP-element group 92: 	56 
    -- CP-element group 92: 	57 
    -- CP-element group 92: 	55 
    -- CP-element group 92: 	52 
    -- CP-element group 92: 	46 
    -- CP-element group 92: 	50 
    -- CP-element group 92:  members (45) 
      -- CP-element group 92: 	 branch_block_stmt_2283/merge_stmt_2552__exit__
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658__entry__
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2640_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2646_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2569_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2599_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2605_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2606_complete/req
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/ptr_deref_2610_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/type_cast_2630_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/addr_of_2637_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_update_start
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2283/assign_stmt_2566_to_assign_stmt_2658/array_obj_ref_2636_final_index_sum_regn_Update/req
      -- CP-element group 92: 	 branch_block_stmt_2283/merge_stmt_2552_PhiAck/$exit
      -- CP-element group 92: 	 branch_block_stmt_2283/merge_stmt_2552_PhiAck/phi_stmt_2553_ack
      -- 
    phi_stmt_2553_ack_7623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2553_ack_0, ack => convTransposeC_CP_6511_elements(92)); -- 
    rr_7383_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7383_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2646_inst_req_0); -- 
    cr_7374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => ptr_deref_2640_store_0_req_1); -- 
    req_7324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => addr_of_2637_final_reg_req_1); -- 
    cr_7388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2646_inst_req_1); -- 
    rr_7149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2569_inst_req_0); -- 
    cr_7154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2569_inst_req_1); -- 
    cr_7168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2599_inst_req_1); -- 
    req_7199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => array_obj_ref_2605_index_offset_req_1); -- 
    req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => addr_of_2606_final_reg_req_1); -- 
    cr_7259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => ptr_deref_2610_load_0_req_1); -- 
    cr_7278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => type_cast_2630_inst_req_1); -- 
    req_7309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_7309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeC_CP_6511_elements(92), ack => array_obj_ref_2636_index_offset_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2512_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2533_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2593_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2624_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2361_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2361_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom62_2635_resized : std_logic_vector(13 downto 0);
    signal R_idxprom62_2635_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_2604_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_2604_scaled : std_logic_vector(13 downto 0);
    signal add18_2575 : std_logic_vector(31 downto 0);
    signal add26_2473 : std_logic_vector(31 downto 0);
    signal add37_2488 : std_logic_vector(31 downto 0);
    signal add52_2545 : std_logic_vector(31 downto 0);
    signal add54_2580 : std_logic_vector(31 downto 0);
    signal add67_2653 : std_logic_vector(31 downto 0);
    signal add_2458 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2605_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2605_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2605_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2605_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2605_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2605_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2636_root_address : std_logic_vector(13 downto 0);
    signal arrayidx63_2638 : std_logic_vector(31 downto 0);
    signal arrayidx_2607 : std_logic_vector(31 downto 0);
    signal call_2286 : std_logic_vector(15 downto 0);
    signal cmp79_2689 : std_logic_vector(0 downto 0);
    signal cmp87_2715 : std_logic_vector(0 downto 0);
    signal cmp_2658 : std_logic_vector(0 downto 0);
    signal conv10100_2570 : std_logic_vector(31 downto 0);
    signal conv13_2443 : std_logic_vector(31 downto 0);
    signal conv16_2448 : std_logic_vector(31 downto 0);
    signal conv23_2347 : std_logic_vector(31 downto 0);
    signal conv28_2366 : std_logic_vector(31 downto 0);
    signal conv34_2380 : std_logic_vector(31 downto 0);
    signal conv47_2514 : std_logic_vector(31 downto 0);
    signal conv50_2535 : std_logic_vector(31 downto 0);
    signal conv66_2647 : std_logic_vector(31 downto 0);
    signal conv76_2684 : std_logic_vector(31 downto 0);
    signal conv85_2710 : std_logic_vector(31 downto 0);
    signal conv_2309 : std_logic_vector(15 downto 0);
    signal div78_2422 : std_logic_vector(31 downto 0);
    signal div_2305 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2412 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2295 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2317 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2329 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2339 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2355 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2372 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2388 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2400 : std_logic_vector(31 downto 0);
    signal idxprom62_2631 : std_logic_vector(63 downto 0);
    signal idxprom_2600 : std_logic_vector(63 downto 0);
    signal inc83_2693 : std_logic_vector(15 downto 0);
    signal inc83x_xinput_dim0x_x2_2698 : std_logic_vector(15 downto 0);
    signal inc_2679 : std_logic_vector(15 downto 0);
    signal indvar_2553 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_2671 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2432 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2425 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_2705 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_2566 : std_logic_vector(15 downto 0);
    signal mul17_2463 : std_logic_vector(31 downto 0);
    signal mul24_2468 : std_logic_vector(31 downto 0);
    signal mul35_2483 : std_logic_vector(31 downto 0);
    signal mul51_2540 : std_logic_vector(31 downto 0);
    signal mul53_2550 : std_logic_vector(31 downto 0);
    signal mul_2453 : std_logic_vector(31 downto 0);
    signal ptr_deref_2298_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2298_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2298_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2298_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2298_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2320_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2320_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2320_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2320_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2320_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2332_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2332_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2332_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2332_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2332_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2342_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2342_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2342_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2342_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2342_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2358_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2358_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2358_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2358_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2358_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2375_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2375_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2375_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2375_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2375_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2391_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2391_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2391_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2391_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2391_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2403_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2403_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2415_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2415_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2415_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2415_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2415_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2610_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2610_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2610_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2610_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2610_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_2640_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_2640_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2640_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext101_2526 : std_logic_vector(31 downto 0);
    signal sext103_2586 : std_logic_vector(31 downto 0);
    signal sext104_2617 : std_logic_vector(31 downto 0);
    signal sext_2505 : std_logic_vector(31 downto 0);
    signal shr61_2626 : std_logic_vector(31 downto 0);
    signal shr_2595 : std_logic_vector(31 downto 0);
    signal sub29_2520 : std_logic_vector(31 downto 0);
    signal sub40_2493 : std_logic_vector(31 downto 0);
    signal sub41_2499 : std_logic_vector(31 downto 0);
    signal sub_2478 : std_logic_vector(31 downto 0);
    signal tmp11_2321 : std_logic_vector(31 downto 0);
    signal tmp14_2333 : std_logic_vector(31 downto 0);
    signal tmp22_2343 : std_logic_vector(15 downto 0);
    signal tmp25_2359 : std_logic_vector(31 downto 0);
    signal tmp27_2362 : std_logic_vector(15 downto 0);
    signal tmp33_2376 : std_logic_vector(15 downto 0);
    signal tmp36_2392 : std_logic_vector(31 downto 0);
    signal tmp45_2404 : std_logic_vector(31 downto 0);
    signal tmp48_2416 : std_logic_vector(31 downto 0);
    signal tmp58_2611 : std_logic_vector(63 downto 0);
    signal tmp_2299 : std_logic_vector(31 downto 0);
    signal type_cast_2303_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2420_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2429_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2431_wire : std_logic_vector(15 downto 0);
    signal type_cast_2435_wire : std_logic_vector(15 downto 0);
    signal type_cast_2437_wire : std_logic_vector(15 downto 0);
    signal type_cast_2441_wire : std_logic_vector(31 downto 0);
    signal type_cast_2446_wire : std_logic_vector(31 downto 0);
    signal type_cast_2497_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2503_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2508_wire : std_logic_vector(31 downto 0);
    signal type_cast_2511_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2518_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2529_wire : std_logic_vector(31 downto 0);
    signal type_cast_2532_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2557_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2559_wire : std_logic_vector(15 downto 0);
    signal type_cast_2564_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2584_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2589_wire : std_logic_vector(31 downto 0);
    signal type_cast_2592_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2598_wire : std_logic_vector(63 downto 0);
    signal type_cast_2615_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2620_wire : std_logic_vector(31 downto 0);
    signal type_cast_2623_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2629_wire : std_logic_vector(63 downto 0);
    signal type_cast_2645_wire : std_logic_vector(31 downto 0);
    signal type_cast_2651_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2669_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2677_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2682_wire : std_logic_vector(31 downto 0);
    signal type_cast_2702_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2708_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2361_word_address_0 <= "0";
    array_obj_ref_2605_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2605_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2605_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2605_resized_base_address <= "00000000000000";
    array_obj_ref_2636_constant_part_of_offset <= "00000000000000";
    array_obj_ref_2636_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_2636_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_2636_resized_base_address <= "00000000000000";
    iNsTr_10_2412 <= "00000000000000000000000000000011";
    iNsTr_2_2295 <= "00000000000000000000000000000010";
    iNsTr_3_2317 <= "00000000000000000000000000000100";
    iNsTr_4_2329 <= "00000000000000000000000000000011";
    iNsTr_5_2339 <= "00000000000000000000000000000000";
    iNsTr_6_2355 <= "00000000000000000000000000000011";
    iNsTr_7_2372 <= "00000000000000000000000000000001";
    iNsTr_8_2388 <= "00000000000000000000000000000100";
    iNsTr_9_2400 <= "00000000000000000000000000000100";
    ptr_deref_2298_word_offset_0 <= "0000000";
    ptr_deref_2320_word_offset_0 <= "0000000";
    ptr_deref_2332_word_offset_0 <= "0000000";
    ptr_deref_2342_word_offset_0 <= "0";
    ptr_deref_2358_word_offset_0 <= "0000000";
    ptr_deref_2375_word_offset_0 <= "0";
    ptr_deref_2391_word_offset_0 <= "0000000";
    ptr_deref_2403_word_offset_0 <= "0000000";
    ptr_deref_2415_word_offset_0 <= "0000000";
    ptr_deref_2610_word_offset_0 <= "00000000000000";
    ptr_deref_2640_word_offset_0 <= "00000000000000";
    type_cast_2303_wire_constant <= "00000000000000000000000000000001";
    type_cast_2420_wire_constant <= "00000000000000000000000000000001";
    type_cast_2429_wire_constant <= "0000000000000000";
    type_cast_2497_wire_constant <= "00000000000000000000000000010000";
    type_cast_2503_wire_constant <= "11111111111111110000000000000000";
    type_cast_2511_wire_constant <= "00000000000000000000000000010000";
    type_cast_2518_wire_constant <= "00000000000000000000000000010000";
    type_cast_2524_wire_constant <= "11111111111111110000000000000000";
    type_cast_2532_wire_constant <= "00000000000000000000000000010000";
    type_cast_2557_wire_constant <= "0000000000000000";
    type_cast_2564_wire_constant <= "0000000000000100";
    type_cast_2584_wire_constant <= "00000000000000000000000000010000";
    type_cast_2592_wire_constant <= "00000000000000000000000000010010";
    type_cast_2615_wire_constant <= "00000000000000000000000000010000";
    type_cast_2623_wire_constant <= "00000000000000000000000000010010";
    type_cast_2651_wire_constant <= "00000000000000000000000000000100";
    type_cast_2669_wire_constant <= "0000000000000001";
    type_cast_2677_wire_constant <= "0000000000000001";
    type_cast_2702_wire_constant <= "0000000000000000";
    phi_stmt_2425: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2429_wire_constant & type_cast_2431_wire;
      req <= phi_stmt_2425_req_0 & phi_stmt_2425_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2425",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2425_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2425,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2425
    phi_stmt_2432: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2435_wire & type_cast_2437_wire;
      req <= phi_stmt_2432_req_0 & phi_stmt_2432_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2432",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2432_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2432,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2432
    phi_stmt_2553: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2557_wire_constant & type_cast_2559_wire;
      req <= phi_stmt_2553_req_0 & phi_stmt_2553_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2553",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2553_ack_0,
          idata => idata,
          odata => indvar_2553,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2553
    -- flow-through select operator MUX_2704_inst
    input_dim1x_x2_2705 <= type_cast_2702_wire_constant when (cmp79_2689(0) /=  '0') else inc_2679;
    addr_of_2606_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2606_final_reg_req_0;
      addr_of_2606_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2606_final_reg_req_1;
      addr_of_2606_final_reg_ack_1<= rack(0);
      addr_of_2606_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2606_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2605_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_2607,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_2637_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_2637_final_reg_req_0;
      addr_of_2637_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_2637_final_reg_req_1;
      addr_of_2637_final_reg_ack_1<= rack(0);
      addr_of_2637_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_2637_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_2636_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx63_2638,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2308_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2308_inst_req_0;
      type_cast_2308_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2308_inst_req_1;
      type_cast_2308_inst_ack_1<= rack(0);
      type_cast_2308_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2308_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2305,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2309,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2346_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2346_inst_req_0;
      type_cast_2346_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2346_inst_req_1;
      type_cast_2346_inst_ack_1<= rack(0);
      type_cast_2346_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2346_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp22_2343,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_2347,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2365_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2365_inst_req_0;
      type_cast_2365_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2365_inst_req_1;
      type_cast_2365_inst_ack_1<= rack(0);
      type_cast_2365_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2365_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp27_2362,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv28_2366,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2379_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2379_inst_req_0;
      type_cast_2379_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2379_inst_req_1;
      type_cast_2379_inst_ack_1<= rack(0);
      type_cast_2379_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2379_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp33_2376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv34_2380,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2431_inst_req_0;
      type_cast_2431_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2431_inst_req_1;
      type_cast_2431_inst_ack_1<= rack(0);
      type_cast_2431_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2431_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_2705,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2431_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2435_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2435_inst_req_0;
      type_cast_2435_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2435_inst_req_1;
      type_cast_2435_inst_ack_1<= rack(0);
      type_cast_2435_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2435_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2435_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2437_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2437_inst_req_0;
      type_cast_2437_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2437_inst_req_1;
      type_cast_2437_inst_ack_1<= rack(0);
      type_cast_2437_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2437_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc83x_xinput_dim0x_x2_2698,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2437_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2442_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2442_inst_req_0;
      type_cast_2442_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2442_inst_req_1;
      type_cast_2442_inst_ack_1<= rack(0);
      type_cast_2442_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2442_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2441_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13_2443,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2447_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2447_inst_req_0;
      type_cast_2447_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2447_inst_req_1;
      type_cast_2447_inst_ack_1<= rack(0);
      type_cast_2447_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2447_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2446_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2448,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2508_inst
    process(sext_2505) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2505(31 downto 0);
      type_cast_2508_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2513_inst
    process(ASHR_i32_i32_2512_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2512_wire(31 downto 0);
      conv47_2514 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2529_inst
    process(sext101_2526) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext101_2526(31 downto 0);
      type_cast_2529_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2534_inst
    process(ASHR_i32_i32_2533_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2533_wire(31 downto 0);
      conv50_2535 <= tmp_var; -- 
    end process;
    type_cast_2559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2559_inst_req_0;
      type_cast_2559_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2559_inst_req_1;
      type_cast_2559_inst_ack_1<= rack(0);
      type_cast_2559_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2559_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_2671,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2559_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2569_inst_req_0;
      type_cast_2569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2569_inst_req_1;
      type_cast_2569_inst_ack_1<= rack(0);
      type_cast_2569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_2566,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv10100_2570,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2589_inst
    process(sext103_2586) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext103_2586(31 downto 0);
      type_cast_2589_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2594_inst
    process(ASHR_i32_i32_2593_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2593_wire(31 downto 0);
      shr_2595 <= tmp_var; -- 
    end process;
    type_cast_2599_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2599_inst_req_0;
      type_cast_2599_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2599_inst_req_1;
      type_cast_2599_inst_ack_1<= rack(0);
      type_cast_2599_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2599_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2598_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_2600,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2620_inst
    process(sext104_2617) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext104_2617(31 downto 0);
      type_cast_2620_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2625_inst
    process(ASHR_i32_i32_2624_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2624_wire(31 downto 0);
      shr61_2626 <= tmp_var; -- 
    end process;
    type_cast_2630_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2630_inst_req_0;
      type_cast_2630_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2630_inst_req_1;
      type_cast_2630_inst_ack_1<= rack(0);
      type_cast_2630_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2630_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2629_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom62_2631,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2646_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2646_inst_req_0;
      type_cast_2646_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2646_inst_req_1;
      type_cast_2646_inst_ack_1<= rack(0);
      type_cast_2646_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2646_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2645_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv66_2647,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2683_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2683_inst_req_0;
      type_cast_2683_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2683_inst_req_1;
      type_cast_2683_inst_ack_1<= rack(0);
      type_cast_2683_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2683_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2682_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv76_2684,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2692_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2692_inst_req_0;
      type_cast_2692_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2692_inst_req_1;
      type_cast_2692_inst_ack_1<= rack(0);
      type_cast_2692_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2692_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => cmp79_2689,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc83_2693,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2709_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2709_inst_req_0;
      type_cast_2709_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2709_inst_req_1;
      type_cast_2709_inst_ack_1<= rack(0);
      type_cast_2709_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2709_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2708_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_2710,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2361_gather_scatter
    process(LOAD_padding_2361_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2361_data_0;
      ov(15 downto 0) := iv;
      tmp27_2362 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2605_index_1_rename
    process(R_idxprom_2604_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_2604_resized;
      ov(13 downto 0) := iv;
      R_idxprom_2604_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2605_index_1_resize
    process(idxprom_2600) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_2600;
      ov := iv(13 downto 0);
      R_idxprom_2604_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2605_root_address_inst
    process(array_obj_ref_2605_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2605_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2605_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_index_1_rename
    process(R_idxprom62_2635_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom62_2635_resized;
      ov(13 downto 0) := iv;
      R_idxprom62_2635_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_index_1_resize
    process(idxprom62_2631) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom62_2631;
      ov := iv(13 downto 0);
      R_idxprom62_2635_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2636_root_address_inst
    process(array_obj_ref_2636_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2636_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_2636_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_addr_0
    process(ptr_deref_2298_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2298_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2298_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_base_resize
    process(iNsTr_2_2295) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2295;
      ov := iv(6 downto 0);
      ptr_deref_2298_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_gather_scatter
    process(ptr_deref_2298_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2298_data_0;
      ov(31 downto 0) := iv;
      tmp_2299 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2298_root_address_inst
    process(ptr_deref_2298_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2298_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2298_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2320_addr_0
    process(ptr_deref_2320_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2320_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2320_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2320_base_resize
    process(iNsTr_3_2317) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2317;
      ov := iv(6 downto 0);
      ptr_deref_2320_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2320_gather_scatter
    process(ptr_deref_2320_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2320_data_0;
      ov(31 downto 0) := iv;
      tmp11_2321 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2320_root_address_inst
    process(ptr_deref_2320_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2320_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2320_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2332_addr_0
    process(ptr_deref_2332_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2332_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2332_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2332_base_resize
    process(iNsTr_4_2329) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2329;
      ov := iv(6 downto 0);
      ptr_deref_2332_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2332_gather_scatter
    process(ptr_deref_2332_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2332_data_0;
      ov(31 downto 0) := iv;
      tmp14_2333 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2332_root_address_inst
    process(ptr_deref_2332_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2332_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2332_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2342_addr_0
    process(ptr_deref_2342_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2342_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2342_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2342_base_resize
    process(iNsTr_5_2339) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2339;
      ov := iv(0 downto 0);
      ptr_deref_2342_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2342_gather_scatter
    process(ptr_deref_2342_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2342_data_0;
      ov(15 downto 0) := iv;
      tmp22_2343 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2342_root_address_inst
    process(ptr_deref_2342_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2342_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2342_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_addr_0
    process(ptr_deref_2358_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2358_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_base_resize
    process(iNsTr_6_2355) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2355;
      ov := iv(6 downto 0);
      ptr_deref_2358_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_gather_scatter
    process(ptr_deref_2358_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_data_0;
      ov(31 downto 0) := iv;
      tmp25_2359 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2358_root_address_inst
    process(ptr_deref_2358_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2358_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2358_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2375_addr_0
    process(ptr_deref_2375_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2375_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2375_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2375_base_resize
    process(iNsTr_7_2372) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2372;
      ov := iv(0 downto 0);
      ptr_deref_2375_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2375_gather_scatter
    process(ptr_deref_2375_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2375_data_0;
      ov(15 downto 0) := iv;
      tmp33_2376 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2375_root_address_inst
    process(ptr_deref_2375_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2375_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2375_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2391_addr_0
    process(ptr_deref_2391_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2391_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2391_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2391_base_resize
    process(iNsTr_8_2388) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2388;
      ov := iv(6 downto 0);
      ptr_deref_2391_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2391_gather_scatter
    process(ptr_deref_2391_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2391_data_0;
      ov(31 downto 0) := iv;
      tmp36_2392 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2391_root_address_inst
    process(ptr_deref_2391_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2391_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2391_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_addr_0
    process(ptr_deref_2403_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2403_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_base_resize
    process(iNsTr_9_2400) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2400;
      ov := iv(6 downto 0);
      ptr_deref_2403_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_gather_scatter
    process(ptr_deref_2403_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_data_0;
      ov(31 downto 0) := iv;
      tmp45_2404 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2403_root_address_inst
    process(ptr_deref_2403_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2403_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2403_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_addr_0
    process(ptr_deref_2415_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2415_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_base_resize
    process(iNsTr_10_2412) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2412;
      ov := iv(6 downto 0);
      ptr_deref_2415_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_gather_scatter
    process(ptr_deref_2415_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_data_0;
      ov(31 downto 0) := iv;
      tmp48_2416 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2415_root_address_inst
    process(ptr_deref_2415_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2415_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2415_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2610_addr_0
    process(ptr_deref_2610_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2610_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2610_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2610_base_resize
    process(arrayidx_2607) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_2607;
      ov := iv(13 downto 0);
      ptr_deref_2610_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2610_gather_scatter
    process(ptr_deref_2610_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2610_data_0;
      ov(63 downto 0) := iv;
      tmp58_2611 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2610_root_address_inst
    process(ptr_deref_2610_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2610_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2610_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_addr_0
    process(ptr_deref_2640_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2640_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_2640_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_base_resize
    process(arrayidx63_2638) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx63_2638;
      ov := iv(13 downto 0);
      ptr_deref_2640_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_gather_scatter
    process(tmp58_2611) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp58_2611;
      ov(63 downto 0) := iv;
      ptr_deref_2640_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2640_root_address_inst
    process(ptr_deref_2640_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2640_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_2640_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_2659_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_2658;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2659_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2659_branch_req_0,
          ack0 => if_stmt_2659_branch_ack_0,
          ack1 => if_stmt_2659_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2716_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp87_2715;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_2716_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2716_branch_req_0,
          ack0 => if_stmt_2716_branch_ack_0,
          ack1 => if_stmt_2716_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_2670_inst
    process(indvar_2553) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_2553, type_cast_2669_wire_constant, tmp_var);
      indvarx_xnext_2671 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2678_inst
    process(input_dim1x_x1x_xph_2425) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2425, type_cast_2677_wire_constant, tmp_var);
      inc_2679 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_2697_inst
    process(inc83_2693, input_dim0x_x2x_xph_2432) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(inc83_2693, input_dim0x_x2x_xph_2432, tmp_var);
      inc83x_xinput_dim0x_x2_2698 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2457_inst
    process(mul_2453, conv13_2443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2453, conv13_2443, tmp_var);
      add_2458 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2472_inst
    process(mul24_2468, tmp25_2359) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul24_2468, tmp25_2359, tmp_var);
      add26_2473 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2487_inst
    process(mul35_2483, tmp36_2392) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul35_2483, tmp36_2392, tmp_var);
      add37_2488 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2504_inst
    process(sub41_2499) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub41_2499, type_cast_2503_wire_constant, tmp_var);
      sext_2505 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2525_inst
    process(sub29_2520) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub29_2520, type_cast_2524_wire_constant, tmp_var);
      sext101_2526 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2544_inst
    process(conv47_2514, mul51_2540) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv47_2514, mul51_2540, tmp_var);
      add52_2545 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2574_inst
    process(mul17_2463, conv10100_2570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul17_2463, conv10100_2570, tmp_var);
      add18_2575 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2579_inst
    process(mul53_2550, conv10100_2570) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul53_2550, conv10100_2570, tmp_var);
      add54_2580 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2652_inst
    process(conv66_2647) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv66_2647, type_cast_2651_wire_constant, tmp_var);
      add67_2653 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2512_inst
    process(type_cast_2508_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2508_wire, type_cast_2511_wire_constant, tmp_var);
      ASHR_i32_i32_2512_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2533_inst
    process(type_cast_2529_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2529_wire, type_cast_2532_wire_constant, tmp_var);
      ASHR_i32_i32_2533_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2593_inst
    process(type_cast_2589_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2589_wire, type_cast_2592_wire_constant, tmp_var);
      ASHR_i32_i32_2593_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2624_inst
    process(type_cast_2620_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2620_wire, type_cast_2623_wire_constant, tmp_var);
      ASHR_i32_i32_2624_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2688_inst
    process(conv76_2684, div78_2422) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv76_2684, div78_2422, tmp_var);
      cmp79_2689 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_2714_inst
    process(conv85_2710, tmp_2299) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv85_2710, tmp_2299, tmp_var);
      cmp87_2715 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2304_inst
    process(tmp_2299) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2299, type_cast_2303_wire_constant, tmp_var);
      div_2305 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2421_inst
    process(tmp14_2333) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp14_2333, type_cast_2420_wire_constant, tmp_var);
      div78_2422 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_2565_inst
    process(indvar_2553) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_2553, type_cast_2564_wire_constant, tmp_var);
      input_dim2x_x1_2566 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2452_inst
    process(tmp14_2333, conv16_2448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp14_2333, conv16_2448, tmp_var);
      mul_2453 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2462_inst
    process(add_2458, tmp11_2321) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2458, tmp11_2321, tmp_var);
      mul17_2463 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2467_inst
    process(conv23_2347, conv16_2448) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv23_2347, conv16_2448, tmp_var);
      mul24_2468 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2482_inst
    process(conv34_2380, conv13_2443) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv34_2380, conv13_2443, tmp_var);
      mul35_2483 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2539_inst
    process(tmp48_2416, conv50_2535) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_2416, conv50_2535, tmp_var);
      mul51_2540 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2549_inst
    process(add52_2545, tmp45_2404) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add52_2545, tmp45_2404, tmp_var);
      mul53_2550 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2498_inst
    process(sub40_2493) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub40_2493, type_cast_2497_wire_constant, tmp_var);
      sub41_2499 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2519_inst
    process(sub_2478) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2478, type_cast_2518_wire_constant, tmp_var);
      sub29_2520 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2585_inst
    process(add18_2575) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add18_2575, type_cast_2584_wire_constant, tmp_var);
      sext103_2586 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2616_inst
    process(add54_2580) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add54_2580, type_cast_2615_wire_constant, tmp_var);
      sext104_2617 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2477_inst
    process(add26_2473, conv28_2366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add26_2473, conv28_2366, tmp_var);
      sub_2478 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2492_inst
    process(add37_2488, conv28_2366) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add37_2488, conv28_2366, tmp_var);
      sub40_2493 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_2657_inst
    process(add67_2653, tmp11_2321) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add67_2653, tmp11_2321, tmp_var);
      cmp_2658 <= tmp_var; --
    end process;
    -- shared split operator group (34) : array_obj_ref_2605_index_offset 
    ApIntAdd_group_34: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_2604_scaled;
      array_obj_ref_2605_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2605_index_offset_req_0;
      array_obj_ref_2605_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2605_index_offset_req_1;
      array_obj_ref_2605_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_34_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_34_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_34",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : array_obj_ref_2636_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom62_2635_scaled;
      array_obj_ref_2636_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_2636_index_offset_req_0;
      array_obj_ref_2636_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_2636_index_offset_req_1;
      array_obj_ref_2636_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- unary operator type_cast_2441_inst
    process(input_dim1x_x1x_xph_2425) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2425, tmp_var);
      type_cast_2441_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2446_inst
    process(input_dim0x_x2x_xph_2432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2432, tmp_var);
      type_cast_2446_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2598_inst
    process(shr_2595) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_2595, tmp_var);
      type_cast_2598_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2629_inst
    process(shr61_2626) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr61_2626, tmp_var);
      type_cast_2629_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2645_inst
    process(input_dim2x_x1_2566) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_2566, tmp_var);
      type_cast_2645_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2682_inst
    process(inc_2679) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_2679, tmp_var);
      type_cast_2682_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2708_inst
    process(inc83x_xinput_dim0x_x2_2698) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc83x_xinput_dim0x_x2_2698, tmp_var);
      type_cast_2708_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2361_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2361_load_0_req_0;
      LOAD_padding_2361_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2361_load_0_req_1;
      LOAD_padding_2361_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2361_word_address_0;
      LOAD_padding_2361_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2298_load_0 ptr_deref_2320_load_0 ptr_deref_2332_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2298_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2320_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2332_load_0_req_0;
      ptr_deref_2298_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2320_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2332_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2298_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2320_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2332_load_0_req_1;
      ptr_deref_2298_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2320_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2332_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2298_word_address_0 & ptr_deref_2320_word_address_0 & ptr_deref_2332_word_address_0;
      ptr_deref_2298_data_0 <= data_out(95 downto 64);
      ptr_deref_2320_data_0 <= data_out(63 downto 32);
      ptr_deref_2332_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2342_load_0 ptr_deref_2375_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2342_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2375_load_0_req_0;
      ptr_deref_2342_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2375_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2342_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2375_load_0_req_1;
      ptr_deref_2342_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2375_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2342_word_address_0 & ptr_deref_2375_word_address_0;
      ptr_deref_2342_data_0 <= data_out(31 downto 16);
      ptr_deref_2375_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2358_load_0 ptr_deref_2391_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2358_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2391_load_0_req_0;
      ptr_deref_2358_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2391_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2358_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2391_load_0_req_1;
      ptr_deref_2358_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2391_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2358_word_address_0 & ptr_deref_2391_word_address_0;
      ptr_deref_2358_data_0 <= data_out(63 downto 32);
      ptr_deref_2391_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2403_load_0 ptr_deref_2415_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2403_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2415_load_0_req_0;
      ptr_deref_2403_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2415_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2403_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2415_load_0_req_1;
      ptr_deref_2403_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2415_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2403_word_address_0 & ptr_deref_2415_word_address_0;
      ptr_deref_2403_data_0 <= data_out(63 downto 32);
      ptr_deref_2415_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2610_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2610_load_0_req_0;
      ptr_deref_2610_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2610_load_0_req_1;
      ptr_deref_2610_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2610_word_address_0;
      ptr_deref_2610_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_2640_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_2640_store_0_req_0;
      ptr_deref_2640_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_2640_store_0_req_1;
      ptr_deref_2640_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_2640_word_address_0;
      data_in <= ptr_deref_2640_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block2_start_2285_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block2_start_2285_inst_req_0;
      RPIPE_Block2_start_2285_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block2_start_2285_inst_req_1;
      RPIPE_Block2_start_2285_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2286 <= data_out(15 downto 0);
      Block2_start_read_0_gI: SplitGuardInterface generic map(name => "Block2_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block2_start_read_0: InputPortRevised -- 
        generic map ( name => "Block2_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block2_start_pipe_read_req(0),
          oack => Block2_start_pipe_read_ack(0),
          odata => Block2_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block2_done_2724_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block2_done_2724_inst_req_0;
      WPIPE_Block2_done_2724_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block2_done_2724_inst_req_1;
      WPIPE_Block2_done_2724_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2286;
      Block2_done_write_0_gI: SplitGuardInterface generic map(name => "Block2_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block2_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block2_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block2_done_pipe_write_req(0),
          oack => Block2_done_pipe_write_ack(0),
          odata => Block2_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeC_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity convTransposeD is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
    memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
    Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
    Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
    Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
    Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
    Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity convTransposeD;
architecture convTransposeD_arch of convTransposeD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal convTransposeD_CP_7664_start: Boolean;
  signal convTransposeD_CP_7664_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal ptr_deref_2850_load_0_req_0 : boolean;
  signal ptr_deref_2862_load_0_ack_1 : boolean;
  signal LOAD_padding_2820_load_0_req_1 : boolean;
  signal ptr_deref_2862_load_0_req_1 : boolean;
  signal ptr_deref_2834_load_0_ack_0 : boolean;
  signal ptr_deref_2834_load_0_req_0 : boolean;
  signal LOAD_padding_2820_load_0_ack_1 : boolean;
  signal type_cast_2805_inst_ack_1 : boolean;
  signal type_cast_2805_inst_req_1 : boolean;
  signal ptr_deref_2817_load_0_ack_1 : boolean;
  signal type_cast_2894_inst_req_1 : boolean;
  signal type_cast_2894_inst_ack_1 : boolean;
  signal ptr_deref_2874_load_0_req_1 : boolean;
  signal ptr_deref_2874_load_0_ack_1 : boolean;
  signal ptr_deref_2817_load_0_req_1 : boolean;
  signal type_cast_2805_inst_req_0 : boolean;
  signal type_cast_2899_inst_ack_0 : boolean;
  signal type_cast_2899_inst_req_0 : boolean;
  signal type_cast_2899_inst_ack_1 : boolean;
  signal type_cast_3021_inst_req_1 : boolean;
  signal type_cast_2805_inst_ack_0 : boolean;
  signal type_cast_3051_inst_ack_1 : boolean;
  signal type_cast_2838_inst_req_0 : boolean;
  signal ptr_deref_2862_load_0_req_0 : boolean;
  signal type_cast_3021_inst_ack_1 : boolean;
  signal type_cast_3021_inst_req_0 : boolean;
  signal type_cast_3051_inst_req_1 : boolean;
  signal type_cast_2894_inst_req_0 : boolean;
  signal type_cast_3021_inst_ack_0 : boolean;
  signal type_cast_2899_inst_req_1 : boolean;
  signal ptr_deref_2817_load_0_req_0 : boolean;
  signal ptr_deref_2817_load_0_ack_0 : boolean;
  signal LOAD_padding_2820_load_0_ack_0 : boolean;
  signal RPIPE_Block3_start_2734_inst_req_0 : boolean;
  signal RPIPE_Block3_start_2734_inst_ack_0 : boolean;
  signal RPIPE_Block3_start_2734_inst_req_1 : boolean;
  signal RPIPE_Block3_start_2734_inst_ack_1 : boolean;
  signal LOAD_padding_2820_load_0_req_0 : boolean;
  signal ptr_deref_2747_load_0_req_0 : boolean;
  signal ptr_deref_2747_load_0_ack_0 : boolean;
  signal ptr_deref_2747_load_0_req_1 : boolean;
  signal ptr_deref_2747_load_0_ack_1 : boolean;
  signal ptr_deref_2874_load_0_ack_0 : boolean;
  signal type_cast_3051_inst_ack_0 : boolean;
  signal ptr_deref_2874_load_0_req_0 : boolean;
  signal type_cast_2757_inst_req_0 : boolean;
  signal type_cast_2757_inst_ack_0 : boolean;
  signal type_cast_2757_inst_req_1 : boolean;
  signal type_cast_2757_inst_ack_1 : boolean;
  signal ptr_deref_2834_load_0_ack_1 : boolean;
  signal ptr_deref_2769_load_0_req_0 : boolean;
  signal ptr_deref_2769_load_0_ack_0 : boolean;
  signal ptr_deref_2769_load_0_req_1 : boolean;
  signal ptr_deref_2769_load_0_ack_1 : boolean;
  signal type_cast_3051_inst_req_0 : boolean;
  signal type_cast_2894_inst_ack_0 : boolean;
  signal type_cast_2779_inst_req_0 : boolean;
  signal type_cast_2779_inst_ack_0 : boolean;
  signal ptr_deref_2834_load_0_req_1 : boolean;
  signal type_cast_2779_inst_req_1 : boolean;
  signal type_cast_2779_inst_ack_1 : boolean;
  signal ptr_deref_2850_load_0_ack_1 : boolean;
  signal ptr_deref_2850_load_0_req_1 : boolean;
  signal type_cast_2838_inst_ack_1 : boolean;
  signal type_cast_2838_inst_req_1 : boolean;
  signal ptr_deref_2791_load_0_req_0 : boolean;
  signal ptr_deref_2791_load_0_ack_0 : boolean;
  signal ptr_deref_2791_load_0_req_1 : boolean;
  signal ptr_deref_2791_load_0_ack_1 : boolean;
  signal ptr_deref_2850_load_0_ack_0 : boolean;
  signal ptr_deref_2862_load_0_ack_0 : boolean;
  signal type_cast_2824_inst_ack_1 : boolean;
  signal type_cast_2824_inst_req_1 : boolean;
  signal type_cast_2824_inst_ack_0 : boolean;
  signal type_cast_2824_inst_req_0 : boolean;
  signal type_cast_2838_inst_ack_0 : boolean;
  signal ptr_deref_2801_load_0_req_0 : boolean;
  signal ptr_deref_2801_load_0_ack_0 : boolean;
  signal ptr_deref_2801_load_0_req_1 : boolean;
  signal ptr_deref_2801_load_0_ack_1 : boolean;
  signal array_obj_ref_3057_index_offset_req_0 : boolean;
  signal array_obj_ref_3057_index_offset_ack_0 : boolean;
  signal array_obj_ref_3057_index_offset_req_1 : boolean;
  signal array_obj_ref_3057_index_offset_ack_1 : boolean;
  signal addr_of_3058_final_reg_req_0 : boolean;
  signal addr_of_3058_final_reg_ack_0 : boolean;
  signal addr_of_3058_final_reg_req_1 : boolean;
  signal addr_of_3058_final_reg_ack_1 : boolean;
  signal ptr_deref_3062_load_0_req_0 : boolean;
  signal ptr_deref_3062_load_0_ack_0 : boolean;
  signal ptr_deref_3062_load_0_req_1 : boolean;
  signal ptr_deref_3062_load_0_ack_1 : boolean;
  signal type_cast_3082_inst_req_0 : boolean;
  signal type_cast_3082_inst_ack_0 : boolean;
  signal type_cast_3082_inst_req_1 : boolean;
  signal type_cast_3082_inst_ack_1 : boolean;
  signal array_obj_ref_3088_index_offset_req_0 : boolean;
  signal array_obj_ref_3088_index_offset_ack_0 : boolean;
  signal array_obj_ref_3088_index_offset_req_1 : boolean;
  signal array_obj_ref_3088_index_offset_ack_1 : boolean;
  signal addr_of_3089_final_reg_req_0 : boolean;
  signal addr_of_3089_final_reg_ack_0 : boolean;
  signal addr_of_3089_final_reg_req_1 : boolean;
  signal addr_of_3089_final_reg_ack_1 : boolean;
  signal ptr_deref_3092_store_0_req_0 : boolean;
  signal ptr_deref_3092_store_0_ack_0 : boolean;
  signal ptr_deref_3092_store_0_req_1 : boolean;
  signal ptr_deref_3092_store_0_ack_1 : boolean;
  signal type_cast_3098_inst_req_0 : boolean;
  signal type_cast_3098_inst_ack_0 : boolean;
  signal type_cast_3098_inst_req_1 : boolean;
  signal type_cast_3098_inst_ack_1 : boolean;
  signal if_stmt_3111_branch_req_0 : boolean;
  signal if_stmt_3111_branch_ack_1 : boolean;
  signal if_stmt_3111_branch_ack_0 : boolean;
  signal type_cast_3135_inst_req_0 : boolean;
  signal type_cast_3135_inst_ack_0 : boolean;
  signal type_cast_3135_inst_req_1 : boolean;
  signal type_cast_3135_inst_ack_1 : boolean;
  signal if_stmt_3142_branch_req_0 : boolean;
  signal if_stmt_3142_branch_ack_1 : boolean;
  signal if_stmt_3142_branch_ack_0 : boolean;
  signal type_cast_3163_inst_req_0 : boolean;
  signal type_cast_3163_inst_ack_0 : boolean;
  signal type_cast_3163_inst_req_1 : boolean;
  signal type_cast_3163_inst_ack_1 : boolean;
  signal type_cast_3183_inst_req_0 : boolean;
  signal type_cast_3183_inst_ack_0 : boolean;
  signal type_cast_3183_inst_req_1 : boolean;
  signal type_cast_3183_inst_ack_1 : boolean;
  signal if_stmt_3190_branch_req_0 : boolean;
  signal if_stmt_3190_branch_ack_1 : boolean;
  signal if_stmt_3190_branch_ack_0 : boolean;
  signal WPIPE_Block3_done_3198_inst_req_0 : boolean;
  signal WPIPE_Block3_done_3198_inst_ack_0 : boolean;
  signal WPIPE_Block3_done_3198_inst_req_1 : boolean;
  signal WPIPE_Block3_done_3198_inst_ack_1 : boolean;
  signal type_cast_2881_inst_req_0 : boolean;
  signal type_cast_2881_inst_ack_0 : boolean;
  signal type_cast_2881_inst_req_1 : boolean;
  signal type_cast_2881_inst_ack_1 : boolean;
  signal phi_stmt_2878_req_0 : boolean;
  signal type_cast_2887_inst_req_0 : boolean;
  signal type_cast_2887_inst_ack_0 : boolean;
  signal type_cast_2887_inst_req_1 : boolean;
  signal type_cast_2887_inst_ack_1 : boolean;
  signal phi_stmt_2884_req_0 : boolean;
  signal type_cast_2883_inst_req_0 : boolean;
  signal type_cast_2883_inst_ack_0 : boolean;
  signal type_cast_2883_inst_req_1 : boolean;
  signal type_cast_2883_inst_ack_1 : boolean;
  signal phi_stmt_2878_req_1 : boolean;
  signal type_cast_2889_inst_req_0 : boolean;
  signal type_cast_2889_inst_ack_0 : boolean;
  signal type_cast_2889_inst_req_1 : boolean;
  signal type_cast_2889_inst_ack_1 : boolean;
  signal phi_stmt_2884_req_1 : boolean;
  signal phi_stmt_2878_ack_0 : boolean;
  signal phi_stmt_2884_ack_0 : boolean;
  signal type_cast_3011_inst_req_0 : boolean;
  signal type_cast_3011_inst_ack_0 : boolean;
  signal type_cast_3011_inst_req_1 : boolean;
  signal type_cast_3011_inst_ack_1 : boolean;
  signal phi_stmt_3005_req_1 : boolean;
  signal phi_stmt_3005_req_0 : boolean;
  signal phi_stmt_3005_ack_0 : boolean;
  signal type_cast_3172_inst_req_0 : boolean;
  signal type_cast_3172_inst_ack_0 : boolean;
  signal type_cast_3172_inst_req_1 : boolean;
  signal type_cast_3172_inst_ack_1 : boolean;
  signal phi_stmt_3167_req_1 : boolean;
  signal type_cast_3178_inst_req_0 : boolean;
  signal type_cast_3178_inst_ack_0 : boolean;
  signal type_cast_3178_inst_req_1 : boolean;
  signal type_cast_3178_inst_ack_1 : boolean;
  signal phi_stmt_3173_req_1 : boolean;
  signal type_cast_3170_inst_req_0 : boolean;
  signal type_cast_3170_inst_ack_0 : boolean;
  signal type_cast_3170_inst_req_1 : boolean;
  signal type_cast_3170_inst_ack_1 : boolean;
  signal phi_stmt_3167_req_0 : boolean;
  signal type_cast_3176_inst_req_0 : boolean;
  signal type_cast_3176_inst_ack_0 : boolean;
  signal type_cast_3176_inst_req_1 : boolean;
  signal type_cast_3176_inst_ack_1 : boolean;
  signal phi_stmt_3173_req_0 : boolean;
  signal phi_stmt_3167_ack_0 : boolean;
  signal phi_stmt_3173_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "convTransposeD_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  convTransposeD_CP_7664_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "convTransposeD_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= convTransposeD_CP_7664_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  convTransposeD_CP_7664: Block -- control-path 
    signal convTransposeD_CP_7664_elements: BooleanArray(116 downto 0);
    -- 
  begin -- 
    convTransposeD_CP_7664_elements(0) <= convTransposeD_CP_7664_start;
    convTransposeD_CP_7664_symbol <= convTransposeD_CP_7664_elements(74);
    -- CP-element group 0:  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2732/branch_block_stmt_2732__entry__
      -- CP-element group 0: 	 branch_block_stmt_2732/assign_stmt_2735__entry__
      -- CP-element group 0: 	 branch_block_stmt_2732/$entry
      -- CP-element group 0: 	 branch_block_stmt_2732/assign_stmt_2735/$entry
      -- CP-element group 0: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Sample/rr
      -- 
    rr_7722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(0), ack => RPIPE_Block3_start_2734_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_update_start_
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Update/cr
      -- 
    ra_7723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2734_inst_ack_0, ack => convTransposeD_CP_7664_elements(1)); -- 
    cr_7727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(1), ack => RPIPE_Block3_start_2734_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	16 
    -- CP-element group 2: 	28 
    -- CP-element group 2: 	26 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	19 
    -- CP-element group 2: 	27 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	12 
    -- CP-element group 2: 	32 
    -- CP-element group 2: 	31 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	30 
    -- CP-element group 2: 	29 
    -- CP-element group 2: 	22 
    -- CP-element group 2: 	17 
    -- CP-element group 2: 	23 
    -- CP-element group 2: 	24 
    -- CP-element group 2: 	20 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	4 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	7 
    -- CP-element group 2: 	8 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	11 
    -- CP-element group 2:  members (268) 
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2735__exit__
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875__entry__
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2735/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2735/RPIPE_Block3_start_2734_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/word_0/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_update_start_
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Update/cr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_word_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_root_address_calculated
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_plus_offset/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_plus_offset/sum_rename_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_base_plus_offset/sum_rename_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_plus_offset/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_addr_resize/base_resize_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_word_addrgen/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_word_addrgen/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_word_addrgen/root_register_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_word_addrgen/root_register_ack
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_addr_resize/base_resize_req
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_addr_resize/$exit
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_addr_resize/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_base_address_resized
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/word_0/rr
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/word_0/$entry
      -- CP-element group 2: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/word_0/cr
      -- 
    ca_7728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_Block3_start_2734_inst_ack_1, ack => convTransposeD_CP_7664_elements(2)); -- 
    rr_8167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2850_load_0_req_0); -- 
    cr_8050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => LOAD_padding_2820_load_0_req_1); -- 
    cr_8228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2862_load_0_req_1); -- 
    rr_8103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2834_load_0_req_0); -- 
    cr_7972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2805_inst_req_1); -- 
    cr_8278_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8278_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2874_load_0_req_1); -- 
    cr_8017_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8017_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2817_load_0_req_1); -- 
    rr_8217_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8217_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2862_load_0_req_0); -- 
    rr_8006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2817_load_0_req_0); -- 
    rr_8039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => LOAD_padding_2820_load_0_req_0); -- 
    rr_7764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2747_load_0_req_0); -- 
    cr_7775_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7775_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2747_load_0_req_1); -- 
    rr_8267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2874_load_0_req_0); -- 
    cr_7794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2757_inst_req_1); -- 
    rr_7828_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7828_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2769_load_0_req_0); -- 
    cr_7839_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7839_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2769_load_0_req_1); -- 
    cr_8114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2834_load_0_req_1); -- 
    cr_7858_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7858_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2779_inst_req_1); -- 
    cr_8178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2850_load_0_req_1); -- 
    cr_8133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2838_inst_req_1); -- 
    rr_7892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2791_load_0_req_0); -- 
    cr_7903_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7903_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2791_load_0_req_1); -- 
    cr_8069_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8069_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => type_cast_2824_inst_req_1); -- 
    rr_7942_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7942_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2801_load_0_req_0); -- 
    cr_7953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_7953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(2), ack => ptr_deref_2801_load_0_req_1); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Sample/word_access_start/word_0/ra
      -- 
    ra_7765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2747_load_0_ack_0, ack => convTransposeD_CP_7664_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (12) 
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/ptr_deref_2747_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/ptr_deref_2747_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/ptr_deref_2747_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2747_Update/ptr_deref_2747_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_sample_start_
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Sample/rr
      -- 
    ca_7776_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2747_load_0_ack_1, ack => convTransposeD_CP_7664_elements(4)); -- 
    rr_7789_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7789_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(4), ack => type_cast_2757_inst_req_0); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Sample/ra
      -- 
    ra_7790_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2757_inst_ack_0, ack => convTransposeD_CP_7664_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	2 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	33 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2757_Update/ca
      -- 
    ca_7795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2757_inst_ack_1, ack => convTransposeD_CP_7664_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/$exit
      -- CP-element group 7: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Sample/word_access_start/word_0/ra
      -- 
    ra_7829_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2769_load_0_ack_0, ack => convTransposeD_CP_7664_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (12) 
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/$exit
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/word_0/$exit
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/word_access_complete/word_0/ca
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/ptr_deref_2769_Merge/$entry
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/ptr_deref_2769_Merge/$exit
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/ptr_deref_2769_Merge/merge_req
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2769_Update/ptr_deref_2769_Merge/merge_ack
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Sample/rr
      -- 
    ca_7840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2769_load_0_ack_1, ack => convTransposeD_CP_7664_elements(8)); -- 
    rr_7853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(8), ack => type_cast_2779_inst_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Sample/ra
      -- 
    ra_7854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2779_inst_ack_0, ack => convTransposeD_CP_7664_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	33 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Update/$exit
      -- CP-element group 10: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2779_Update/ca
      -- 
    ca_7859_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2779_inst_ack_1, ack => convTransposeD_CP_7664_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (5) 
      -- CP-element group 11: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_sample_completed_
      -- CP-element group 11: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/$exit
      -- CP-element group 11: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/$exit
      -- CP-element group 11: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/word_0/$exit
      -- CP-element group 11: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Sample/word_access_start/word_0/ra
      -- 
    ra_7893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2791_load_0_ack_0, ack => convTransposeD_CP_7664_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	2 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	33 
    -- CP-element group 12:  members (9) 
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_update_completed_
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/$exit
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/$exit
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/word_0/$exit
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/word_access_complete/word_0/ca
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/ptr_deref_2791_Merge/$entry
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/ptr_deref_2791_Merge/$exit
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/ptr_deref_2791_Merge/merge_req
      -- CP-element group 12: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2791_Update/ptr_deref_2791_Merge/merge_ack
      -- 
    ca_7904_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2791_load_0_ack_1, ack => convTransposeD_CP_7664_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/$exit
      -- CP-element group 13: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/word_0/$exit
      -- CP-element group 13: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Sample/word_access_start/word_0/ra
      -- 
    ra_7943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2801_load_0_ack_0, ack => convTransposeD_CP_7664_elements(13)); -- 
    -- CP-element group 14:  transition  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (12) 
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/$exit
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/word_0/$exit
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/word_access_complete/word_0/ca
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/ptr_deref_2801_Merge/$entry
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/ptr_deref_2801_Merge/$exit
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/ptr_deref_2801_Merge/merge_req
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2801_Update/ptr_deref_2801_Merge/merge_ack
      -- CP-element group 14: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_sample_start_
      -- 
    ca_7954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2801_load_0_ack_1, ack => convTransposeD_CP_7664_elements(14)); -- 
    rr_7967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_7967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(14), ack => type_cast_2805_inst_req_0); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_sample_completed_
      -- 
    ra_7968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2805_inst_ack_0, ack => convTransposeD_CP_7664_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	2 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	33 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Update/ca
      -- CP-element group 16: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2805_update_completed_
      -- 
    ca_7973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2805_inst_ack_1, ack => convTransposeD_CP_7664_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	2 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (5) 
      -- CP-element group 17: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/word_0/ra
      -- CP-element group 17: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/word_access_start/$exit
      -- CP-element group 17: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Sample/$exit
      -- 
    ra_8007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2817_load_0_ack_0, ack => convTransposeD_CP_7664_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	2 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	33 
    -- CP-element group 18:  members (9) 
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/word_0/ca
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/ptr_deref_2817_Merge/$entry
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/ptr_deref_2817_Merge/$exit
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/ptr_deref_2817_Merge/merge_req
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/ptr_deref_2817_Merge/merge_ack
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/word_0/$exit
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/word_access_complete/$exit
      -- CP-element group 18: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2817_Update/$exit
      -- 
    ca_8018_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2817_load_0_ack_1, ack => convTransposeD_CP_7664_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	2 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (5) 
      -- CP-element group 19: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/word_0/ra
      -- CP-element group 19: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/word_0/$exit
      -- CP-element group 19: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/word_access_start/$exit
      -- CP-element group 19: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Sample/$exit
      -- 
    ra_8040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2820_load_0_ack_0, ack => convTransposeD_CP_7664_elements(19)); -- 
    -- CP-element group 20:  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	2 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (12) 
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/LOAD_padding_2820_Merge/$exit
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/LOAD_padding_2820_Merge/$entry
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/word_0/ca
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/word_0/$exit
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/LOAD_padding_2820_Merge/merge_req
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/word_access_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/LOAD_padding_2820_Merge/merge_ack
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/LOAD_padding_2820_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Sample/rr
      -- CP-element group 20: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Sample/$entry
      -- 
    ca_8051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => LOAD_padding_2820_load_0_ack_1, ack => convTransposeD_CP_7664_elements(20)); -- 
    rr_8064_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8064_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(20), ack => type_cast_2824_inst_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Sample/ra
      -- CP-element group 21: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Sample/$exit
      -- 
    ra_8065_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2824_inst_ack_0, ack => convTransposeD_CP_7664_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	33 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Update/ca
      -- CP-element group 22: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2824_Update/$exit
      -- 
    ca_8070_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2824_inst_ack_1, ack => convTransposeD_CP_7664_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	2 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/word_0/ra
      -- CP-element group 23: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/word_0/$exit
      -- CP-element group 23: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/word_access_start/$exit
      -- CP-element group 23: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_sample_completed_
      -- 
    ra_8104_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_0_ack_0, ack => convTransposeD_CP_7664_elements(23)); -- 
    -- CP-element group 24:  transition  input  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	2 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (12) 
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/$exit
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Sample/rr
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/ptr_deref_2834_Merge/merge_ack
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/ptr_deref_2834_Merge/merge_req
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/ptr_deref_2834_Merge/$exit
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/ptr_deref_2834_Merge/$entry
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/word_0/ca
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_Update/word_access_complete/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2834_update_completed_
      -- 
    ca_8115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_0_ack_1, ack => convTransposeD_CP_7664_elements(24)); -- 
    rr_8128_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8128_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(24), ack => type_cast_2838_inst_req_0); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Sample/ra
      -- 
    ra_8129_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2838_inst_ack_0, ack => convTransposeD_CP_7664_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	2 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	33 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/type_cast_2838_Update/$exit
      -- 
    ca_8134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2838_inst_ack_1, ack => convTransposeD_CP_7664_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	2 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (5) 
      -- CP-element group 27: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/word_0/$exit
      -- CP-element group 27: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/$exit
      -- CP-element group 27: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Sample/word_access_start/word_0/ra
      -- 
    ra_8168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2850_load_0_ack_0, ack => convTransposeD_CP_7664_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	33 
    -- CP-element group 28:  members (9) 
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/ptr_deref_2850_Merge/merge_ack
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/ptr_deref_2850_Merge/merge_req
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/ptr_deref_2850_Merge/$exit
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/ptr_deref_2850_Merge/$entry
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/word_0/ca
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/word_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/word_access_complete/$exit
      -- CP-element group 28: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2850_Update/$exit
      -- 
    ca_8179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2850_load_0_ack_1, ack => convTransposeD_CP_7664_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	2 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/$exit
      -- CP-element group 29: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/word_0/$exit
      -- CP-element group 29: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Sample/word_access_start/word_0/ra
      -- 
    ra_8218_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2862_load_0_ack_0, ack => convTransposeD_CP_7664_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	2 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	33 
    -- CP-element group 30:  members (9) 
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/ptr_deref_2862_Merge/$entry
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/word_0/ca
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/word_0/$exit
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/word_access_complete/$exit
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/ptr_deref_2862_Merge/merge_ack
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/ptr_deref_2862_Merge/merge_req
      -- CP-element group 30: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2862_Update/ptr_deref_2862_Merge/$exit
      -- 
    ca_8229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2862_load_0_ack_1, ack => convTransposeD_CP_7664_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/word_0/ra
      -- CP-element group 31: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Sample/$exit
      -- 
    ra_8268_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2874_load_0_ack_0, ack => convTransposeD_CP_7664_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	2 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	33 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/ptr_deref_2874_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/ptr_deref_2874_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/ptr_deref_2874_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_Update/ptr_deref_2874_Merge/merge_ack
      -- CP-element group 32: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/ptr_deref_2874_update_completed_
      -- 
    ca_8279_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2874_load_0_ack_1, ack => convTransposeD_CP_7664_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  place  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	16 
    -- CP-element group 33: 	28 
    -- CP-element group 33: 	26 
    -- CP-element group 33: 	18 
    -- CP-element group 33: 	12 
    -- CP-element group 33: 	32 
    -- CP-element group 33: 	30 
    -- CP-element group 33: 	22 
    -- CP-element group 33: 	6 
    -- CP-element group 33: 	10 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	75 
    -- CP-element group 33: 	76 
    -- CP-element group 33: 	78 
    -- CP-element group 33: 	79 
    -- CP-element group 33:  members (20) 
      -- CP-element group 33: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875__exit__
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter
      -- CP-element group 33: 	 branch_block_stmt_2732/assign_stmt_2744_to_assign_stmt_2875/$exit
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Update/cr
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Update/cr
      -- 
    rr_8713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2881_inst_req_0); -- 
    cr_8718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2881_inst_req_1); -- 
    rr_8736_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8736_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2887_inst_req_0); -- 
    cr_8741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(33), ack => type_cast_2887_inst_req_1); -- 
    convTransposeD_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(16) & convTransposeD_CP_7664_elements(28) & convTransposeD_CP_7664_elements(26) & convTransposeD_CP_7664_elements(18) & convTransposeD_CP_7664_elements(12) & convTransposeD_CP_7664_elements(32) & convTransposeD_CP_7664_elements(30) & convTransposeD_CP_7664_elements(22) & convTransposeD_CP_7664_elements(6) & convTransposeD_CP_7664_elements(10);
      gj_convTransposeD_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	92 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Sample/ra
      -- 
    ra_8296_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2894_inst_ack_0, ack => convTransposeD_CP_7664_elements(34)); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	92 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	38 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Update/ca
      -- CP-element group 35: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Update/$exit
      -- 
    ca_8301_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2894_inst_ack_1, ack => convTransposeD_CP_7664_elements(35)); -- 
    -- CP-element group 36:  transition  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	92 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_sample_completed_
      -- CP-element group 36: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Sample/ra
      -- 
    ra_8310_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2899_inst_ack_0, ack => convTransposeD_CP_7664_elements(36)); -- 
    -- CP-element group 37:  transition  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	92 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_update_completed_
      -- CP-element group 37: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Update/ca
      -- CP-element group 37: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Update/$exit
      -- 
    ca_8315_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2899_inst_ack_1, ack => convTransposeD_CP_7664_elements(37)); -- 
    -- CP-element group 38:  join  transition  place  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	35 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	96 
    -- CP-element group 38:  members (6) 
      -- CP-element group 38: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/$exit
      -- CP-element group 38: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody
      -- CP-element group 38: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002__exit__
      -- CP-element group 38: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$entry
      -- CP-element group 38: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/$entry
      -- CP-element group 38: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$entry
      -- 
    convTransposeD_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(35) & convTransposeD_CP_7664_elements(37);
      gj_convTransposeD_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	98 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Sample/ra
      -- 
    ra_8327_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3021_inst_ack_0, ack => convTransposeD_CP_7664_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	98 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40: 	49 
    -- CP-element group 40:  members (9) 
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Update/ca
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Sample/rr
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Sample/rr
      -- 
    ca_8332_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3021_inst_ack_1, ack => convTransposeD_CP_7664_elements(40)); -- 
    rr_8340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(40), ack => type_cast_3051_inst_req_0); -- 
    rr_8450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(40), ack => type_cast_3082_inst_req_0); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Sample/ra
      -- 
    ra_8341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_0, ack => convTransposeD_CP_7664_elements(41)); -- 
    -- CP-element group 42:  transition  input  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	98 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (16) 
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Update/ca
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_resized_1
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_scaled_1
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_computed_1
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_resize_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_resize_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_resize_1/index_resize_req
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_resize_1/index_resize_ack
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_scale_1/$entry
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_scale_1/$exit
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_scale_1/scale_rename_req
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_index_scale_1/scale_rename_ack
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Sample/req
      -- 
    ca_8346_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3051_inst_ack_1, ack => convTransposeD_CP_7664_elements(42)); -- 
    req_8371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(42), ack => array_obj_ref_3057_index_offset_req_0); -- 
    -- CP-element group 43:  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	60 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_sample_complete
      -- CP-element group 43: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Sample/ack
      -- 
    ack_8372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3057_index_offset_ack_0, ack => convTransposeD_CP_7664_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	98 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (11) 
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_root_address_calculated
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_offset_calculated
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Update/ack
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_base_plus_offset/$entry
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_base_plus_offset/$exit
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_base_plus_offset/sum_rename_req
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_base_plus_offset/sum_rename_ack
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_request/$entry
      -- CP-element group 44: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_request/req
      -- 
    ack_8377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3057_index_offset_ack_1, ack => convTransposeD_CP_7664_elements(44)); -- 
    req_8386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(44), ack => addr_of_3058_final_reg_req_0); -- 
    -- CP-element group 45:  transition  input  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_request/$exit
      -- CP-element group 45: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_request/ack
      -- 
    ack_8387_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3058_final_reg_ack_0, ack => convTransposeD_CP_7664_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	98 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (24) 
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_update_completed_
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_complete/$exit
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_complete/ack
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_word_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_root_address_calculated
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_address_resized
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_addr_resize/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_addr_resize/$exit
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_addr_resize/base_resize_req
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_addr_resize/base_resize_ack
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_plus_offset/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_plus_offset/$exit
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_plus_offset/sum_rename_req
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_base_plus_offset/sum_rename_ack
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_word_addrgen/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_word_addrgen/$exit
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_word_addrgen/root_register_req
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_word_addrgen/root_register_ack
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/word_0/$entry
      -- CP-element group 46: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/word_0/rr
      -- 
    ack_8392_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3058_final_reg_ack_1, ack => convTransposeD_CP_7664_elements(46)); -- 
    rr_8425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(46), ack => ptr_deref_3062_load_0_req_0); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (5) 
      -- CP-element group 47: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/$exit
      -- CP-element group 47: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/word_0/$exit
      -- CP-element group 47: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Sample/word_access_start/word_0/ra
      -- 
    ra_8426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3062_load_0_ack_0, ack => convTransposeD_CP_7664_elements(47)); -- 
    -- CP-element group 48:  transition  input  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	98 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	55 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/$exit
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/word_0/$exit
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/word_0/ca
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/ptr_deref_3062_Merge/$entry
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/ptr_deref_3062_Merge/$exit
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/ptr_deref_3062_Merge/merge_req
      -- CP-element group 48: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/ptr_deref_3062_Merge/merge_ack
      -- 
    ca_8437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3062_load_0_ack_1, ack => convTransposeD_CP_7664_elements(48)); -- 
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	40 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Sample/ra
      -- 
    ra_8451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3082_inst_ack_0, ack => convTransposeD_CP_7664_elements(49)); -- 
    -- CP-element group 50:  transition  input  output  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	98 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (16) 
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Update/ca
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_resized_1
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_scaled_1
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_computed_1
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_resize_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_resize_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_resize_1/index_resize_req
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_resize_1/index_resize_ack
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_scale_1/$entry
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_scale_1/$exit
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_scale_1/scale_rename_req
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_index_scale_1/scale_rename_ack
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Sample/req
      -- 
    ca_8456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3082_inst_ack_1, ack => convTransposeD_CP_7664_elements(50)); -- 
    req_8481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(50), ack => array_obj_ref_3088_index_offset_req_0); -- 
    -- CP-element group 51:  transition  input  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	60 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_sample_complete
      -- CP-element group 51: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Sample/ack
      -- 
    ack_8482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3088_index_offset_ack_0, ack => convTransposeD_CP_7664_elements(51)); -- 
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	98 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (11) 
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_request/$entry
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_root_address_calculated
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_offset_calculated
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_base_plus_offset/$entry
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_base_plus_offset/$exit
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_base_plus_offset/sum_rename_req
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_base_plus_offset/sum_rename_ack
      -- CP-element group 52: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_request/req
      -- 
    ack_8487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3088_index_offset_ack_1, ack => convTransposeD_CP_7664_elements(52)); -- 
    req_8496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(52), ack => addr_of_3089_final_reg_req_0); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_request/$exit
      -- CP-element group 53: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_request/ack
      -- 
    ack_8497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3089_final_reg_ack_0, ack => convTransposeD_CP_7664_elements(53)); -- 
    -- CP-element group 54:  fork  transition  input  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	98 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (19) 
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_complete/$exit
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_complete/ack
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_word_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_root_address_calculated
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_address_resized
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_addr_resize/$entry
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_addr_resize/$exit
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_addr_resize/base_resize_req
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_addr_resize/base_resize_ack
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_plus_offset/$entry
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_plus_offset/$exit
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_plus_offset/sum_rename_req
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_base_plus_offset/sum_rename_ack
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_word_addrgen/$entry
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_word_addrgen/$exit
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_word_addrgen/root_register_req
      -- CP-element group 54: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_word_addrgen/root_register_ack
      -- 
    ack_8502_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3089_final_reg_ack_1, ack => convTransposeD_CP_7664_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	48 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (9) 
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/ptr_deref_3092_Split/$entry
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/ptr_deref_3092_Split/$exit
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/ptr_deref_3092_Split/split_req
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/ptr_deref_3092_Split/split_ack
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/$entry
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/word_0/$entry
      -- CP-element group 55: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/word_0/rr
      -- 
    rr_8540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(55), ack => ptr_deref_3092_store_0_req_0); -- 
    convTransposeD_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(48) & convTransposeD_CP_7664_elements(54);
      gj_convTransposeD_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (5) 
      -- CP-element group 56: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/$exit
      -- CP-element group 56: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/word_0/$exit
      -- CP-element group 56: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Sample/word_access_start/word_0/ra
      -- 
    ra_8541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3092_store_0_ack_0, ack => convTransposeD_CP_7664_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	98 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	60 
    -- CP-element group 57:  members (5) 
      -- CP-element group 57: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/$exit
      -- CP-element group 57: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/word_0/$exit
      -- CP-element group 57: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/word_0/ca
      -- 
    ca_8552_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3092_store_0_ack_1, ack => convTransposeD_CP_7664_elements(57)); -- 
    -- CP-element group 58:  transition  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	98 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Sample/ra
      -- 
    ra_8561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3098_inst_ack_0, ack => convTransposeD_CP_7664_elements(58)); -- 
    -- CP-element group 59:  transition  input  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	98 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Update/ca
      -- 
    ca_8566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3098_inst_ack_1, ack => convTransposeD_CP_7664_elements(59)); -- 
    -- CP-element group 60:  branch  join  transition  place  output  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	43 
    -- CP-element group 60: 	51 
    -- CP-element group 60: 	57 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (10) 
      -- CP-element group 60: 	 branch_block_stmt_2732/R_cmp_3112_place
      -- CP-element group 60: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/$exit
      -- CP-element group 60: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110__exit__
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111__entry__
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_dead_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_eval_test/$entry
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_eval_test/$exit
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_eval_test/branch_req
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_if_link/$entry
      -- CP-element group 60: 	 branch_block_stmt_2732/if_stmt_3111_else_link/$entry
      -- 
    branch_req_8574_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8574_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(60), ack => if_stmt_3111_branch_req_0); -- 
    convTransposeD_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(43) & convTransposeD_CP_7664_elements(51) & convTransposeD_CP_7664_elements(57) & convTransposeD_CP_7664_elements(59);
      gj_convTransposeD_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	94 
    -- CP-element group 61: 	93 
    -- CP-element group 61:  members (24) 
      -- CP-element group 61: 	 branch_block_stmt_2732/whilex_xbody_ifx_xthen
      -- CP-element group 61: 	 branch_block_stmt_2732/merge_stmt_3117__exit__
      -- CP-element group 61: 	 branch_block_stmt_2732/assign_stmt_3123__entry__
      -- CP-element group 61: 	 branch_block_stmt_2732/assign_stmt_3123__exit__
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody
      -- CP-element group 61: 	 branch_block_stmt_2732/if_stmt_3111_if_link/$exit
      -- CP-element group 61: 	 branch_block_stmt_2732/if_stmt_3111_if_link/if_choice_transition
      -- CP-element group 61: 	 branch_block_stmt_2732/assign_stmt_3123/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/assign_stmt_3123/$exit
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Update/cr
      -- CP-element group 61: 	 branch_block_stmt_2732/whilex_xbody_ifx_xthen_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/whilex_xbody_ifx_xthen_PhiReq/$exit
      -- CP-element group 61: 	 branch_block_stmt_2732/merge_stmt_3117_PhiReqMerge
      -- CP-element group 61: 	 branch_block_stmt_2732/merge_stmt_3117_PhiAck/$entry
      -- CP-element group 61: 	 branch_block_stmt_2732/merge_stmt_3117_PhiAck/$exit
      -- CP-element group 61: 	 branch_block_stmt_2732/merge_stmt_3117_PhiAck/dummy
      -- 
    if_choice_transition_8579_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3111_branch_ack_1, ack => convTransposeD_CP_7664_elements(61)); -- 
    rr_8817_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8817_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(61), ack => type_cast_3011_inst_req_0); -- 
    cr_8822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(61), ack => type_cast_3011_inst_req_1); -- 
    -- CP-element group 62:  fork  transition  place  input  output  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (18) 
      -- CP-element group 62: 	 branch_block_stmt_2732/merge_stmt_3125__exit__
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141__entry__
      -- CP-element group 62: 	 branch_block_stmt_2732/if_stmt_3111_else_link/$exit
      -- CP-element group 62: 	 branch_block_stmt_2732/if_stmt_3111_else_link/else_choice_transition
      -- CP-element group 62: 	 branch_block_stmt_2732/whilex_xbody_ifx_xelse
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/$entry
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_update_start_
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Sample/rr
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Update/$entry
      -- CP-element group 62: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_2732/whilex_xbody_ifx_xelse_PhiReq/$entry
      -- CP-element group 62: 	 branch_block_stmt_2732/whilex_xbody_ifx_xelse_PhiReq/$exit
      -- CP-element group 62: 	 branch_block_stmt_2732/merge_stmt_3125_PhiReqMerge
      -- CP-element group 62: 	 branch_block_stmt_2732/merge_stmt_3125_PhiAck/$entry
      -- CP-element group 62: 	 branch_block_stmt_2732/merge_stmt_3125_PhiAck/$exit
      -- CP-element group 62: 	 branch_block_stmt_2732/merge_stmt_3125_PhiAck/dummy
      -- 
    else_choice_transition_8583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3111_branch_ack_0, ack => convTransposeD_CP_7664_elements(62)); -- 
    rr_8599_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8599_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(62), ack => type_cast_3135_inst_req_0); -- 
    cr_8604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(62), ack => type_cast_3135_inst_req_1); -- 
    -- CP-element group 63:  transition  input  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Sample/ra
      -- 
    ra_8600_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3135_inst_ack_0, ack => convTransposeD_CP_7664_elements(63)); -- 
    -- CP-element group 64:  branch  transition  place  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (13) 
      -- CP-element group 64: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141__exit__
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142__entry__
      -- CP-element group 64: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/$exit
      -- CP-element group 64: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Update/$exit
      -- CP-element group 64: 	 branch_block_stmt_2732/assign_stmt_3131_to_assign_stmt_3141/type_cast_3135_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_dead_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_eval_test/$entry
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_eval_test/$exit
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_eval_test/branch_req
      -- CP-element group 64: 	 branch_block_stmt_2732/R_cmp81_3143_place
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_if_link/$entry
      -- CP-element group 64: 	 branch_block_stmt_2732/if_stmt_3142_else_link/$entry
      -- 
    ca_8605_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3135_inst_ack_1, ack => convTransposeD_CP_7664_elements(64)); -- 
    branch_req_8613_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8613_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(64), ack => if_stmt_3142_branch_req_0); -- 
    -- CP-element group 65:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: 	68 
    -- CP-element group 65:  members (18) 
      -- CP-element group 65: 	 branch_block_stmt_2732/merge_stmt_3148__exit__
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164__entry__
      -- CP-element group 65: 	 branch_block_stmt_2732/if_stmt_3142_if_link/$exit
      -- CP-element group 65: 	 branch_block_stmt_2732/if_stmt_3142_if_link/if_choice_transition
      -- CP-element group 65: 	 branch_block_stmt_2732/ifx_xelse_ifx_xthen83
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/$entry
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_update_start_
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Sample/rr
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_2732/ifx_xelse_ifx_xthen83_PhiReq/$entry
      -- CP-element group 65: 	 branch_block_stmt_2732/ifx_xelse_ifx_xthen83_PhiReq/$exit
      -- CP-element group 65: 	 branch_block_stmt_2732/merge_stmt_3148_PhiReqMerge
      -- CP-element group 65: 	 branch_block_stmt_2732/merge_stmt_3148_PhiAck/$entry
      -- CP-element group 65: 	 branch_block_stmt_2732/merge_stmt_3148_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_2732/merge_stmt_3148_PhiAck/dummy
      -- 
    if_choice_transition_8618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3142_branch_ack_1, ack => convTransposeD_CP_7664_elements(65)); -- 
    rr_8635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(65), ack => type_cast_3163_inst_req_0); -- 
    cr_8640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(65), ack => type_cast_3163_inst_req_1); -- 
    -- CP-element group 66:  fork  transition  place  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	99 
    -- CP-element group 66: 	100 
    -- CP-element group 66: 	102 
    -- CP-element group 66: 	103 
    -- CP-element group 66:  members (20) 
      -- CP-element group 66: 	 branch_block_stmt_2732/if_stmt_3142_else_link/$exit
      -- CP-element group 66: 	 branch_block_stmt_2732/if_stmt_3142_else_link/else_choice_transition
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Update/cr
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Sample/rr
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3142_branch_ack_0, ack => convTransposeD_CP_7664_elements(66)); -- 
    rr_8891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3172_inst_req_0); -- 
    cr_8896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3172_inst_req_1); -- 
    rr_8914_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8914_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3178_inst_req_0); -- 
    cr_8919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(66), ack => type_cast_3178_inst_req_1); -- 
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Sample/ra
      -- 
    ra_8636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3163_inst_ack_0, ack => convTransposeD_CP_7664_elements(67)); -- 
    -- CP-element group 68:  fork  transition  place  input  output  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	65 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	109 
    -- CP-element group 68: 	110 
    -- CP-element group 68: 	107 
    -- CP-element group 68: 	106 
    -- CP-element group 68:  members (23) 
      -- CP-element group 68: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164__exit__
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend
      -- CP-element group 68: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/$exit
      -- CP-element group 68: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2732/assign_stmt_3154_to_assign_stmt_3164/type_cast_3163_Update/ca
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Update/cr
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Sample/rr
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Update/cr
      -- 
    ca_8641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3163_inst_ack_1, ack => convTransposeD_CP_7664_elements(68)); -- 
    rr_8940_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8940_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3170_inst_req_0); -- 
    cr_8945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3170_inst_req_1); -- 
    rr_8963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3176_inst_req_0); -- 
    cr_8968_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8968_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(68), ack => type_cast_3176_inst_req_1); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	116 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_sample_completed_
      -- CP-element group 69: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Sample/$exit
      -- CP-element group 69: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Sample/ra
      -- 
    ra_8653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_0, ack => convTransposeD_CP_7664_elements(69)); -- 
    -- CP-element group 70:  branch  transition  place  input  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	116 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (13) 
      -- CP-element group 70: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189__exit__
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190__entry__
      -- CP-element group 70: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/$exit
      -- CP-element group 70: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_update_completed_
      -- CP-element group 70: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Update/$exit
      -- CP-element group 70: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Update/ca
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_2732/R_cmp92_3191_place
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_2732/if_stmt_3190_else_link/$entry
      -- 
    ca_8658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3183_inst_ack_1, ack => convTransposeD_CP_7664_elements(70)); -- 
    branch_req_8666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_8666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(70), ack => if_stmt_3190_branch_req_0); -- 
    -- CP-element group 71:  merge  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (15) 
      -- CP-element group 71: 	 branch_block_stmt_2732/merge_stmt_3196__exit__
      -- CP-element group 71: 	 branch_block_stmt_2732/assign_stmt_3200__entry__
      -- CP-element group 71: 	 branch_block_stmt_2732/if_stmt_3190_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_2732/if_stmt_3190_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_2732/ifx_xend_whilex_xend
      -- CP-element group 71: 	 branch_block_stmt_2732/assign_stmt_3200/$entry
      -- CP-element group 71: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_sample_start_
      -- CP-element group 71: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Sample/req
      -- CP-element group 71: 	 branch_block_stmt_2732/ifx_xend_whilex_xend_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_2732/ifx_xend_whilex_xend_PhiReq/$exit
      -- CP-element group 71: 	 branch_block_stmt_2732/merge_stmt_3196_PhiReqMerge
      -- CP-element group 71: 	 branch_block_stmt_2732/merge_stmt_3196_PhiAck/$entry
      -- CP-element group 71: 	 branch_block_stmt_2732/merge_stmt_3196_PhiAck/$exit
      -- CP-element group 71: 	 branch_block_stmt_2732/merge_stmt_3196_PhiAck/dummy
      -- 
    if_choice_transition_8671_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3190_branch_ack_1, ack => convTransposeD_CP_7664_elements(71)); -- 
    req_8688_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8688_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(71), ack => WPIPE_Block3_done_3198_inst_req_0); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	82 
    -- CP-element group 72: 	83 
    -- CP-element group 72: 	85 
    -- CP-element group 72: 	86 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_2732/if_stmt_3190_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_2732/if_stmt_3190_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Update/cr
      -- 
    else_choice_transition_8675_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3190_branch_ack_0, ack => convTransposeD_CP_7664_elements(72)); -- 
    rr_8762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2883_inst_req_0); -- 
    cr_8767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2883_inst_req_1); -- 
    rr_8785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2889_inst_req_0); -- 
    cr_8790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(72), ack => type_cast_2889_inst_req_1); -- 
    -- CP-element group 73:  transition  input  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (6) 
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_sample_completed_
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_update_start_
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Sample/$exit
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Sample/ack
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Update/req
      -- 
    ack_8689_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3198_inst_ack_0, ack => convTransposeD_CP_7664_elements(73)); -- 
    req_8693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(73), ack => WPIPE_Block3_done_3198_inst_req_1); -- 
    -- CP-element group 74:  transition  place  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (16) 
      -- CP-element group 74: 	 $exit
      -- CP-element group 74: 	 branch_block_stmt_2732/branch_block_stmt_2732__exit__
      -- CP-element group 74: 	 branch_block_stmt_2732/$exit
      -- CP-element group 74: 	 branch_block_stmt_2732/assign_stmt_3200__exit__
      -- CP-element group 74: 	 branch_block_stmt_2732/return__
      -- CP-element group 74: 	 branch_block_stmt_2732/merge_stmt_3202__exit__
      -- CP-element group 74: 	 branch_block_stmt_2732/assign_stmt_3200/$exit
      -- CP-element group 74: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_update_completed_
      -- CP-element group 74: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Update/$exit
      -- CP-element group 74: 	 branch_block_stmt_2732/assign_stmt_3200/WPIPE_Block3_done_3198_Update/ack
      -- CP-element group 74: 	 branch_block_stmt_2732/return___PhiReq/$entry
      -- CP-element group 74: 	 branch_block_stmt_2732/return___PhiReq/$exit
      -- CP-element group 74: 	 branch_block_stmt_2732/merge_stmt_3202_PhiReqMerge
      -- CP-element group 74: 	 branch_block_stmt_2732/merge_stmt_3202_PhiAck/$entry
      -- CP-element group 74: 	 branch_block_stmt_2732/merge_stmt_3202_PhiAck/$exit
      -- CP-element group 74: 	 branch_block_stmt_2732/merge_stmt_3202_PhiAck/dummy
      -- 
    ack_8694_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_Block3_done_3198_inst_ack_1, ack => convTransposeD_CP_7664_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	33 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Sample/ra
      -- 
    ra_8714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2881_inst_ack_0, ack => convTransposeD_CP_7664_elements(75)); -- 
    -- CP-element group 76:  transition  input  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	33 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (2) 
      -- CP-element group 76: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/Update/ca
      -- 
    ca_8719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2881_inst_ack_1, ack => convTransposeD_CP_7664_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	81 
    -- CP-element group 77:  members (5) 
      -- CP-element group 77: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/$exit
      -- CP-element group 77: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/$exit
      -- CP-element group 77: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/$exit
      -- CP-element group 77: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2881/SplitProtocol/$exit
      -- CP-element group 77: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_req
      -- 
    phi_stmt_2878_req_8720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2878_req_8720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(77), ack => phi_stmt_2878_req_0); -- 
    convTransposeD_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(75) & convTransposeD_CP_7664_elements(76);
      gj_convTransposeD_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	33 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Sample/ra
      -- 
    ra_8737_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2887_inst_ack_0, ack => convTransposeD_CP_7664_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	33 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/Update/ca
      -- 
    ca_8742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2887_inst_ack_1, ack => convTransposeD_CP_7664_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (5) 
      -- CP-element group 80: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/$exit
      -- CP-element group 80: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/$exit
      -- CP-element group 80: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/$exit
      -- CP-element group 80: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2887/SplitProtocol/$exit
      -- CP-element group 80: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_req
      -- 
    phi_stmt_2884_req_8743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2884_req_8743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(80), ack => phi_stmt_2884_req_0); -- 
    convTransposeD_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(78) & convTransposeD_CP_7664_elements(79);
      gj_convTransposeD_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	77 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	89 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2732/entry_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(77) & convTransposeD_CP_7664_elements(80);
      gj_convTransposeD_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	72 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Sample/ra
      -- 
    ra_8763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2883_inst_ack_0, ack => convTransposeD_CP_7664_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	72 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/Update/ca
      -- 
    ca_8768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2883_inst_ack_1, ack => convTransposeD_CP_7664_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	88 
    -- CP-element group 84:  members (5) 
      -- CP-element group 84: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/$exit
      -- CP-element group 84: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/$exit
      -- CP-element group 84: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/$exit
      -- CP-element group 84: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_sources/type_cast_2883/SplitProtocol/$exit
      -- CP-element group 84: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2878/phi_stmt_2878_req
      -- 
    phi_stmt_2878_req_8769_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2878_req_8769_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(84), ack => phi_stmt_2878_req_1); -- 
    convTransposeD_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(82) & convTransposeD_CP_7664_elements(83);
      gj_convTransposeD_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	72 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Sample/ra
      -- 
    ra_8786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2889_inst_ack_0, ack => convTransposeD_CP_7664_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	72 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (2) 
      -- CP-element group 86: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/Update/ca
      -- 
    ca_8791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2889_inst_ack_1, ack => convTransposeD_CP_7664_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	86 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (5) 
      -- CP-element group 87: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/$exit
      -- CP-element group 87: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/$exit
      -- CP-element group 87: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/$exit
      -- CP-element group 87: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_sources/type_cast_2889/SplitProtocol/$exit
      -- CP-element group 87: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/phi_stmt_2884/phi_stmt_2884_req
      -- 
    phi_stmt_2884_req_8792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2884_req_8792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(87), ack => phi_stmt_2884_req_1); -- 
    convTransposeD_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(85) & convTransposeD_CP_7664_elements(86);
      gj_convTransposeD_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	84 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	89 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2732/ifx_xend_whilex_xbodyx_xouter_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(84) & convTransposeD_CP_7664_elements(87);
      gj_convTransposeD_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  merge  fork  transition  place  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	81 
    -- CP-element group 89: 	88 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	90 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_2732/merge_stmt_2877_PhiReqMerge
      -- CP-element group 89: 	 branch_block_stmt_2732/merge_stmt_2877_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(89) <= OrReduce(convTransposeD_CP_7664_elements(81) & convTransposeD_CP_7664_elements(88));
    -- CP-element group 90:  transition  input  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	89 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_2732/merge_stmt_2877_PhiAck/phi_stmt_2878_ack
      -- 
    phi_stmt_2878_ack_8797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2878_ack_0, ack => convTransposeD_CP_7664_elements(90)); -- 
    -- CP-element group 91:  transition  input  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (1) 
      -- CP-element group 91: 	 branch_block_stmt_2732/merge_stmt_2877_PhiAck/phi_stmt_2884_ack
      -- 
    phi_stmt_2884_ack_8798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2884_ack_0, ack => convTransposeD_CP_7664_elements(91)); -- 
    -- CP-element group 92:  join  fork  transition  place  output  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	34 
    -- CP-element group 92: 	35 
    -- CP-element group 92: 	36 
    -- CP-element group 92: 	37 
    -- CP-element group 92:  members (16) 
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/$entry
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_update_start_
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002__entry__
      -- CP-element group 92: 	 branch_block_stmt_2732/merge_stmt_2877__exit__
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Sample/rr
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2899_Update/cr
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_2732/assign_stmt_2895_to_assign_stmt_3002/type_cast_2894_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_2732/merge_stmt_2877_PhiAck/$exit
      -- 
    cr_8300_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8300_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2894_inst_req_1); -- 
    rr_8309_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8309_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2899_inst_req_0); -- 
    rr_8295_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8295_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2894_inst_req_0); -- 
    cr_8314_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8314_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(92), ack => type_cast_2899_inst_req_1); -- 
    convTransposeD_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(90) & convTransposeD_CP_7664_elements(91);
      gj_convTransposeD_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	61 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (2) 
      -- CP-element group 93: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Sample/ra
      -- 
    ra_8818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_0, ack => convTransposeD_CP_7664_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	61 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (2) 
      -- CP-element group 94: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/Update/ca
      -- 
    ca_8823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3011_inst_ack_1, ack => convTransposeD_CP_7664_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (6) 
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/$exit
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/$exit
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$exit
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/$exit
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3011/SplitProtocol/$exit
      -- CP-element group 95: 	 branch_block_stmt_2732/ifx_xthen_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_req
      -- 
    phi_stmt_3005_req_8824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3005_req_8824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(95), ack => phi_stmt_3005_req_1); -- 
    convTransposeD_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "convTransposeD_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(94) & convTransposeD_CP_7664_elements(93);
      gj_convTransposeD_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  transition  output  delay-element  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	38 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	97 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/$exit
      -- CP-element group 96: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/$exit
      -- CP-element group 96: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/$exit
      -- CP-element group 96: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_sources/type_cast_3009_konst_delay_trans
      -- CP-element group 96: 	 branch_block_stmt_2732/whilex_xbodyx_xouter_whilex_xbody_PhiReq/phi_stmt_3005/phi_stmt_3005_req
      -- 
    phi_stmt_3005_req_8835_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3005_req_8835_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(96), ack => phi_stmt_3005_req_0); -- 
    -- Element group convTransposeD_CP_7664_elements(96) is a control-delay.
    cp_element_96_delay: control_delay_element  generic map(name => " 96_delay", delay_value => 1)  port map(req => convTransposeD_CP_7664_elements(38), ack => convTransposeD_CP_7664_elements(96), clk => clk, reset =>reset);
    -- CP-element group 97:  merge  transition  place  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	96 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	98 
    -- CP-element group 97:  members (2) 
      -- CP-element group 97: 	 branch_block_stmt_2732/merge_stmt_3004_PhiReqMerge
      -- CP-element group 97: 	 branch_block_stmt_2732/merge_stmt_3004_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(97) <= OrReduce(convTransposeD_CP_7664_elements(95) & convTransposeD_CP_7664_elements(96));
    -- CP-element group 98:  fork  transition  place  input  output  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	97 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	50 
    -- CP-element group 98: 	46 
    -- CP-element group 98: 	48 
    -- CP-element group 98: 	42 
    -- CP-element group 98: 	52 
    -- CP-element group 98: 	54 
    -- CP-element group 98: 	57 
    -- CP-element group 98: 	58 
    -- CP-element group 98: 	59 
    -- CP-element group 98: 	39 
    -- CP-element group 98: 	40 
    -- CP-element group 98: 	44 
    -- CP-element group 98:  members (45) 
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/merge_stmt_3004__exit__
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110__entry__
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3021_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3051_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3057_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3058_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3062_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3082_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_update_start
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/array_obj_ref_3088_final_index_sum_regn_Update/req
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/addr_of_3089_complete/req
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/word_0/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/ptr_deref_3092_Update/word_access_complete/word_0/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_sample_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_update_start_
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Sample/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Sample/rr
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Update/$entry
      -- CP-element group 98: 	 branch_block_stmt_2732/assign_stmt_3018_to_assign_stmt_3110/type_cast_3098_Update/cr
      -- CP-element group 98: 	 branch_block_stmt_2732/merge_stmt_3004_PhiAck/$exit
      -- CP-element group 98: 	 branch_block_stmt_2732/merge_stmt_3004_PhiAck/phi_stmt_3005_ack
      -- 
    phi_stmt_3005_ack_8840_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3005_ack_0, ack => convTransposeD_CP_7664_elements(98)); -- 
    cr_8331_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8331_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3021_inst_req_1); -- 
    rr_8326_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8326_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3021_inst_req_0); -- 
    cr_8345_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8345_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3051_inst_req_1); -- 
    req_8376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => array_obj_ref_3057_index_offset_req_1); -- 
    req_8391_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8391_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => addr_of_3058_final_reg_req_1); -- 
    cr_8436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => ptr_deref_3062_load_0_req_1); -- 
    cr_8455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3082_inst_req_1); -- 
    req_8486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => array_obj_ref_3088_index_offset_req_1); -- 
    req_8501_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_8501_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => addr_of_3089_final_reg_req_1); -- 
    cr_8551_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8551_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => ptr_deref_3092_store_0_req_1); -- 
    rr_8560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3098_inst_req_0); -- 
    cr_8565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(98), ack => type_cast_3098_inst_req_1); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	66 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Sample/ra
      -- 
    ra_8892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3172_inst_ack_0, ack => convTransposeD_CP_7664_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	66 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100:  members (2) 
      -- CP-element group 100: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Update/$exit
      -- CP-element group 100: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/Update/ca
      -- 
    ca_8897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3172_inst_ack_1, ack => convTransposeD_CP_7664_elements(100)); -- 
    -- CP-element group 101:  join  transition  output  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	105 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/$exit
      -- CP-element group 101: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/$exit
      -- CP-element group 101: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/$exit
      -- CP-element group 101: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3172/SplitProtocol/$exit
      -- CP-element group 101: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_req
      -- 
    phi_stmt_3167_req_8898_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3167_req_8898_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(101), ack => phi_stmt_3167_req_1); -- 
    convTransposeD_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(99) & convTransposeD_CP_7664_elements(100);
      gj_convTransposeD_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	66 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Sample/$exit
      -- CP-element group 102: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Sample/ra
      -- 
    ra_8915_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3178_inst_ack_0, ack => convTransposeD_CP_7664_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	66 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Update/$exit
      -- CP-element group 103: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/Update/ca
      -- 
    ca_8920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3178_inst_ack_1, ack => convTransposeD_CP_7664_elements(103)); -- 
    -- CP-element group 104:  join  transition  output  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	105 
    -- CP-element group 104:  members (5) 
      -- CP-element group 104: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/$exit
      -- CP-element group 104: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/$exit
      -- CP-element group 104: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/$exit
      -- CP-element group 104: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3178/SplitProtocol/$exit
      -- CP-element group 104: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_req
      -- 
    phi_stmt_3173_req_8921_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3173_req_8921_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(104), ack => phi_stmt_3173_req_1); -- 
    convTransposeD_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(102) & convTransposeD_CP_7664_elements(103);
      gj_convTransposeD_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  join  transition  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	101 
    -- CP-element group 105: 	104 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	113 
    -- CP-element group 105:  members (1) 
      -- CP-element group 105: 	 branch_block_stmt_2732/ifx_xelse_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_105: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_105"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(101) & convTransposeD_CP_7664_elements(104);
      gj_convTransposeD_cp_element_group_105 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(105), clk => clk, reset => reset); --
    end block;
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	68 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Sample/$exit
      -- CP-element group 106: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Sample/ra
      -- 
    ra_8941_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3170_inst_ack_0, ack => convTransposeD_CP_7664_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	68 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	108 
    -- CP-element group 107:  members (2) 
      -- CP-element group 107: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/Update/ca
      -- 
    ca_8946_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3170_inst_ack_1, ack => convTransposeD_CP_7664_elements(107)); -- 
    -- CP-element group 108:  join  transition  output  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	107 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	112 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/$exit
      -- CP-element group 108: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/$exit
      -- CP-element group 108: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/$exit
      -- CP-element group 108: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_sources/type_cast_3170/SplitProtocol/$exit
      -- CP-element group 108: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3167/phi_stmt_3167_req
      -- 
    phi_stmt_3167_req_8947_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3167_req_8947_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(108), ack => phi_stmt_3167_req_0); -- 
    convTransposeD_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(107) & convTransposeD_CP_7664_elements(106);
      gj_convTransposeD_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	68 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (2) 
      -- CP-element group 109: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Sample/ra
      -- 
    ra_8964_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3176_inst_ack_0, ack => convTransposeD_CP_7664_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	68 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	111 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/Update/ca
      -- 
    ca_8969_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3176_inst_ack_1, ack => convTransposeD_CP_7664_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: 	110 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	112 
    -- CP-element group 111:  members (5) 
      -- CP-element group 111: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/$exit
      -- CP-element group 111: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/$exit
      -- CP-element group 111: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/$exit
      -- CP-element group 111: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_sources/type_cast_3176/SplitProtocol/$exit
      -- CP-element group 111: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/phi_stmt_3173/phi_stmt_3173_req
      -- 
    phi_stmt_3173_req_8970_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3173_req_8970_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(111), ack => phi_stmt_3173_req_0); -- 
    convTransposeD_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(109) & convTransposeD_CP_7664_elements(110);
      gj_convTransposeD_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	111 
    -- CP-element group 112: 	108 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	113 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2732/ifx_xthen83_ifx_xend_PhiReq/$exit
      -- 
    convTransposeD_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(111) & convTransposeD_CP_7664_elements(108);
      gj_convTransposeD_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  merge  fork  transition  place  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	112 
    -- CP-element group 113: 	105 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113: 	115 
    -- CP-element group 113:  members (2) 
      -- CP-element group 113: 	 branch_block_stmt_2732/merge_stmt_3166_PhiReqMerge
      -- CP-element group 113: 	 branch_block_stmt_2732/merge_stmt_3166_PhiAck/$entry
      -- 
    convTransposeD_CP_7664_elements(113) <= OrReduce(convTransposeD_CP_7664_elements(112) & convTransposeD_CP_7664_elements(105));
    -- CP-element group 114:  transition  input  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	116 
    -- CP-element group 114:  members (1) 
      -- CP-element group 114: 	 branch_block_stmt_2732/merge_stmt_3166_PhiAck/phi_stmt_3167_ack
      -- 
    phi_stmt_3167_ack_8975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3167_ack_0, ack => convTransposeD_CP_7664_elements(114)); -- 
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	113 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115:  members (1) 
      -- CP-element group 115: 	 branch_block_stmt_2732/merge_stmt_3166_PhiAck/phi_stmt_3173_ack
      -- 
    phi_stmt_3173_ack_8976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3173_ack_0, ack => convTransposeD_CP_7664_elements(115)); -- 
    -- CP-element group 116:  join  fork  transition  place  output  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	114 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	69 
    -- CP-element group 116: 	70 
    -- CP-element group 116:  members (10) 
      -- CP-element group 116: 	 branch_block_stmt_2732/merge_stmt_3166__exit__
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189__entry__
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/$entry
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_sample_start_
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_update_start_
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Sample/$entry
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Sample/rr
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_2732/assign_stmt_3184_to_assign_stmt_3189/type_cast_3183_Update/cr
      -- CP-element group 116: 	 branch_block_stmt_2732/merge_stmt_3166_PhiAck/$exit
      -- 
    rr_8652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_8652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(116), ack => type_cast_3183_inst_req_0); -- 
    cr_8657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_8657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => convTransposeD_CP_7664_elements(116), ack => type_cast_3183_inst_req_1); -- 
    convTransposeD_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "convTransposeD_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= convTransposeD_CP_7664_elements(114) & convTransposeD_CP_7664_elements(115);
      gj_convTransposeD_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => convTransposeD_CP_7664_elements(116), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ASHR_i32_i32_2964_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_2985_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3045_wire : std_logic_vector(31 downto 0);
    signal ASHR_i32_i32_3076_wire : std_logic_vector(31 downto 0);
    signal LOAD_padding_2820_data_0 : std_logic_vector(15 downto 0);
    signal LOAD_padding_2820_word_address_0 : std_logic_vector(0 downto 0);
    signal R_idxprom65_3087_resized : std_logic_vector(13 downto 0);
    signal R_idxprom65_3087_scaled : std_logic_vector(13 downto 0);
    signal R_idxprom_3056_resized : std_logic_vector(13 downto 0);
    signal R_idxprom_3056_scaled : std_logic_vector(13 downto 0);
    signal add21_3027 : std_logic_vector(31 downto 0);
    signal add29_2925 : std_logic_vector(31 downto 0);
    signal add40_2940 : std_logic_vector(31 downto 0);
    signal add55_2997 : std_logic_vector(31 downto 0);
    signal add57_3032 : std_logic_vector(31 downto 0);
    signal add70_3105 : std_logic_vector(31 downto 0);
    signal add_2910 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3057_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3057_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3057_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3057_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3057_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3057_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_3088_root_address : std_logic_vector(13 downto 0);
    signal arrayidx66_3090 : std_logic_vector(31 downto 0);
    signal arrayidx_3059 : std_logic_vector(31 downto 0);
    signal call_2735 : std_logic_vector(15 downto 0);
    signal cmp81_3141 : std_logic_vector(0 downto 0);
    signal cmp92_3189 : std_logic_vector(0 downto 0);
    signal cmp_3110 : std_logic_vector(0 downto 0);
    signal conv13105_3022 : std_logic_vector(31 downto 0);
    signal conv16_2895 : std_logic_vector(31 downto 0);
    signal conv19_2900 : std_logic_vector(31 downto 0);
    signal conv26_2806 : std_logic_vector(31 downto 0);
    signal conv31_2825 : std_logic_vector(31 downto 0);
    signal conv37_2839 : std_logic_vector(31 downto 0);
    signal conv4_2780 : std_logic_vector(15 downto 0);
    signal conv50_2966 : std_logic_vector(31 downto 0);
    signal conv53_2987 : std_logic_vector(31 downto 0);
    signal conv69_3099 : std_logic_vector(31 downto 0);
    signal conv79_3136 : std_logic_vector(31 downto 0);
    signal conv88_3164 : std_logic_vector(15 downto 0);
    signal conv90_3184 : std_logic_vector(31 downto 0);
    signal conv_2758 : std_logic_vector(15 downto 0);
    signal div3_2776 : std_logic_vector(31 downto 0);
    signal div87_3160 : std_logic_vector(31 downto 0);
    signal div_2754 : std_logic_vector(31 downto 0);
    signal iNsTr_10_2871 : std_logic_vector(31 downto 0);
    signal iNsTr_2_2744 : std_logic_vector(31 downto 0);
    signal iNsTr_3_2766 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2788 : std_logic_vector(31 downto 0);
    signal iNsTr_5_2798 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2814 : std_logic_vector(31 downto 0);
    signal iNsTr_7_2831 : std_logic_vector(31 downto 0);
    signal iNsTr_8_2847 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2859 : std_logic_vector(31 downto 0);
    signal idxprom65_3083 : std_logic_vector(63 downto 0);
    signal idxprom_3052 : std_logic_vector(63 downto 0);
    signal inc85_3154 : std_logic_vector(15 downto 0);
    signal inc_3131 : std_logic_vector(15 downto 0);
    signal indvar_3005 : std_logic_vector(15 downto 0);
    signal indvarx_xnext_3123 : std_logic_vector(15 downto 0);
    signal input_dim0x_x0_3173 : std_logic_vector(15 downto 0);
    signal input_dim0x_x2x_xph_2884 : std_logic_vector(15 downto 0);
    signal input_dim1x_x1x_xph_2878 : std_logic_vector(15 downto 0);
    signal input_dim1x_x2_3167 : std_logic_vector(15 downto 0);
    signal input_dim2x_x1_3018 : std_logic_vector(15 downto 0);
    signal mul20_2915 : std_logic_vector(31 downto 0);
    signal mul27_2920 : std_logic_vector(31 downto 0);
    signal mul38_2935 : std_logic_vector(31 downto 0);
    signal mul54_2992 : std_logic_vector(31 downto 0);
    signal mul56_3002 : std_logic_vector(31 downto 0);
    signal mul_2905 : std_logic_vector(31 downto 0);
    signal ptr_deref_2747_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2747_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2747_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2747_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2747_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2769_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2769_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2769_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2769_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2769_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2791_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2791_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2801_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2801_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2801_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2801_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2801_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2817_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2817_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2817_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2817_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2817_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2834_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2834_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_2834_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2834_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_2850_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2850_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2850_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2850_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2850_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2862_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2862_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2862_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2862_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2862_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2874_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2874_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2874_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_2874_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_2874_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_3062_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3062_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3062_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3062_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3062_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_3092_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3092_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_3092_word_offset_0 : std_logic_vector(13 downto 0);
    signal sext106_2978 : std_logic_vector(31 downto 0);
    signal sext108_3038 : std_logic_vector(31 downto 0);
    signal sext109_3069 : std_logic_vector(31 downto 0);
    signal sext_2957 : std_logic_vector(31 downto 0);
    signal shr64_3078 : std_logic_vector(31 downto 0);
    signal shr_3047 : std_logic_vector(31 downto 0);
    signal sub32_2972 : std_logic_vector(31 downto 0);
    signal sub43_2945 : std_logic_vector(31 downto 0);
    signal sub44_2951 : std_logic_vector(31 downto 0);
    signal sub_2930 : std_logic_vector(31 downto 0);
    signal tmp14_2792 : std_logic_vector(31 downto 0);
    signal tmp25_2802 : std_logic_vector(15 downto 0);
    signal tmp28_2818 : std_logic_vector(31 downto 0);
    signal tmp2_2770 : std_logic_vector(31 downto 0);
    signal tmp30_2821 : std_logic_vector(15 downto 0);
    signal tmp36_2835 : std_logic_vector(15 downto 0);
    signal tmp39_2851 : std_logic_vector(31 downto 0);
    signal tmp48_2863 : std_logic_vector(31 downto 0);
    signal tmp51_2875 : std_logic_vector(31 downto 0);
    signal tmp61_3063 : std_logic_vector(63 downto 0);
    signal tmp_2748 : std_logic_vector(31 downto 0);
    signal type_cast_2752_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2774_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2881_wire : std_logic_vector(15 downto 0);
    signal type_cast_2883_wire : std_logic_vector(15 downto 0);
    signal type_cast_2887_wire : std_logic_vector(15 downto 0);
    signal type_cast_2889_wire : std_logic_vector(15 downto 0);
    signal type_cast_2893_wire : std_logic_vector(31 downto 0);
    signal type_cast_2898_wire : std_logic_vector(31 downto 0);
    signal type_cast_2949_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2955_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2960_wire : std_logic_vector(31 downto 0);
    signal type_cast_2963_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2970_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2976_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2981_wire : std_logic_vector(31 downto 0);
    signal type_cast_2984_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3009_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3011_wire : std_logic_vector(15 downto 0);
    signal type_cast_3016_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3036_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3041_wire : std_logic_vector(31 downto 0);
    signal type_cast_3044_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3050_wire : std_logic_vector(63 downto 0);
    signal type_cast_3067_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3072_wire : std_logic_vector(31 downto 0);
    signal type_cast_3075_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3081_wire : std_logic_vector(63 downto 0);
    signal type_cast_3097_wire : std_logic_vector(31 downto 0);
    signal type_cast_3103_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3121_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3129_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3134_wire : std_logic_vector(31 downto 0);
    signal type_cast_3152_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3158_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3170_wire : std_logic_vector(15 downto 0);
    signal type_cast_3172_wire : std_logic_vector(15 downto 0);
    signal type_cast_3176_wire : std_logic_vector(15 downto 0);
    signal type_cast_3178_wire : std_logic_vector(15 downto 0);
    signal type_cast_3182_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    LOAD_padding_2820_word_address_0 <= "0";
    array_obj_ref_3057_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3057_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3057_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3057_resized_base_address <= "00000000000000";
    array_obj_ref_3088_constant_part_of_offset <= "00000000000000";
    array_obj_ref_3088_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_3088_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_3088_resized_base_address <= "00000000000000";
    iNsTr_10_2871 <= "00000000000000000000000000000011";
    iNsTr_2_2744 <= "00000000000000000000000000000010";
    iNsTr_3_2766 <= "00000000000000000000000000000011";
    iNsTr_4_2788 <= "00000000000000000000000000000100";
    iNsTr_5_2798 <= "00000000000000000000000000000000";
    iNsTr_6_2814 <= "00000000000000000000000000000011";
    iNsTr_7_2831 <= "00000000000000000000000000000001";
    iNsTr_8_2847 <= "00000000000000000000000000000100";
    iNsTr_9_2859 <= "00000000000000000000000000000100";
    ptr_deref_2747_word_offset_0 <= "0000000";
    ptr_deref_2769_word_offset_0 <= "0000000";
    ptr_deref_2791_word_offset_0 <= "0000000";
    ptr_deref_2801_word_offset_0 <= "0";
    ptr_deref_2817_word_offset_0 <= "0000000";
    ptr_deref_2834_word_offset_0 <= "0";
    ptr_deref_2850_word_offset_0 <= "0000000";
    ptr_deref_2862_word_offset_0 <= "0000000";
    ptr_deref_2874_word_offset_0 <= "0000000";
    ptr_deref_3062_word_offset_0 <= "00000000000000";
    ptr_deref_3092_word_offset_0 <= "00000000000000";
    type_cast_2752_wire_constant <= "00000000000000000000000000000001";
    type_cast_2774_wire_constant <= "00000000000000000000000000000001";
    type_cast_2949_wire_constant <= "00000000000000000000000000010000";
    type_cast_2955_wire_constant <= "11111111111111110000000000000000";
    type_cast_2963_wire_constant <= "00000000000000000000000000010000";
    type_cast_2970_wire_constant <= "00000000000000000000000000010000";
    type_cast_2976_wire_constant <= "11111111111111110000000000000000";
    type_cast_2984_wire_constant <= "00000000000000000000000000010000";
    type_cast_3009_wire_constant <= "0000000000000000";
    type_cast_3016_wire_constant <= "0000000000000100";
    type_cast_3036_wire_constant <= "00000000000000000000000000010000";
    type_cast_3044_wire_constant <= "00000000000000000000000000010010";
    type_cast_3067_wire_constant <= "00000000000000000000000000010000";
    type_cast_3075_wire_constant <= "00000000000000000000000000010010";
    type_cast_3103_wire_constant <= "00000000000000000000000000000100";
    type_cast_3121_wire_constant <= "0000000000000001";
    type_cast_3129_wire_constant <= "0000000000000001";
    type_cast_3152_wire_constant <= "0000000000000001";
    type_cast_3158_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_2878: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2881_wire & type_cast_2883_wire;
      req <= phi_stmt_2878_req_0 & phi_stmt_2878_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2878",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2878_ack_0,
          idata => idata,
          odata => input_dim1x_x1x_xph_2878,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2878
    phi_stmt_2884: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2887_wire & type_cast_2889_wire;
      req <= phi_stmt_2884_req_0 & phi_stmt_2884_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2884",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2884_ack_0,
          idata => idata,
          odata => input_dim0x_x2x_xph_2884,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2884
    phi_stmt_3005: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3009_wire_constant & type_cast_3011_wire;
      req <= phi_stmt_3005_req_0 & phi_stmt_3005_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3005",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3005_ack_0,
          idata => idata,
          odata => indvar_3005,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3005
    phi_stmt_3167: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3170_wire & type_cast_3172_wire;
      req <= phi_stmt_3167_req_0 & phi_stmt_3167_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3167",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3167_ack_0,
          idata => idata,
          odata => input_dim1x_x2_3167,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3167
    phi_stmt_3173: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3176_wire & type_cast_3178_wire;
      req <= phi_stmt_3173_req_0 & phi_stmt_3173_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3173",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3173_ack_0,
          idata => idata,
          odata => input_dim0x_x0_3173,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3173
    addr_of_3058_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3058_final_reg_req_0;
      addr_of_3058_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3058_final_reg_req_1;
      addr_of_3058_final_reg_ack_1<= rack(0);
      addr_of_3058_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3058_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3057_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_3059,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_3089_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_3089_final_reg_req_0;
      addr_of_3089_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_3089_final_reg_req_1;
      addr_of_3089_final_reg_ack_1<= rack(0);
      addr_of_3089_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_3089_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_3088_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx66_3090,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2757_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2757_inst_req_0;
      type_cast_2757_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2757_inst_req_1;
      type_cast_2757_inst_ack_1<= rack(0);
      type_cast_2757_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2757_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div_2754,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_2758,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2779_inst_req_0;
      type_cast_2779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2779_inst_req_1;
      type_cast_2779_inst_ack_1<= rack(0);
      type_cast_2779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div3_2776,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_2780,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2805_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2805_inst_req_0;
      type_cast_2805_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2805_inst_req_1;
      type_cast_2805_inst_ack_1<= rack(0);
      type_cast_2805_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2805_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp25_2802,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv26_2806,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2824_inst_req_0;
      type_cast_2824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2824_inst_req_1;
      type_cast_2824_inst_ack_1<= rack(0);
      type_cast_2824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp30_2821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv31_2825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2838_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2838_inst_req_0;
      type_cast_2838_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2838_inst_req_1;
      type_cast_2838_inst_ack_1<= rack(0);
      type_cast_2838_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2838_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp36_2835,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv37_2839,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2881_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2881_inst_req_0;
      type_cast_2881_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2881_inst_req_1;
      type_cast_2881_inst_ack_1<= rack(0);
      type_cast_2881_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2881_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_2780,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2881_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2883_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2883_inst_req_0;
      type_cast_2883_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2883_inst_req_1;
      type_cast_2883_inst_ack_1<= rack(0);
      type_cast_2883_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2883_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim1x_x2_3167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2883_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2887_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2887_inst_req_0;
      type_cast_2887_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2887_inst_req_1;
      type_cast_2887_inst_ack_1<= rack(0);
      type_cast_2887_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2887_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv_2758,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2887_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2889_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2889_inst_req_0;
      type_cast_2889_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2889_inst_req_1;
      type_cast_2889_inst_ack_1<= rack(0);
      type_cast_2889_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2889_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x0_3173,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_2889_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2894_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2894_inst_req_0;
      type_cast_2894_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2894_inst_req_1;
      type_cast_2894_inst_ack_1<= rack(0);
      type_cast_2894_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2894_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2893_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_2895,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_2899_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_2899_inst_req_0;
      type_cast_2899_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_2899_inst_req_1;
      type_cast_2899_inst_ack_1<= rack(0);
      type_cast_2899_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_2899_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_2898_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv19_2900,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_2960_inst
    process(sext_2957) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext_2957(31 downto 0);
      type_cast_2960_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2965_inst
    process(ASHR_i32_i32_2964_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2964_wire(31 downto 0);
      conv50_2966 <= tmp_var; -- 
    end process;
    -- interlock type_cast_2981_inst
    process(sext106_2978) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext106_2978(31 downto 0);
      type_cast_2981_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_2986_inst
    process(ASHR_i32_i32_2985_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_2985_wire(31 downto 0);
      conv53_2987 <= tmp_var; -- 
    end process;
    type_cast_3011_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3011_inst_req_0;
      type_cast_3011_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3011_inst_req_1;
      type_cast_3011_inst_ack_1<= rack(0);
      type_cast_3011_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3011_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_3123,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3011_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3021_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3021_inst_req_0;
      type_cast_3021_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3021_inst_req_1;
      type_cast_3021_inst_ack_1<= rack(0);
      type_cast_3021_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3021_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim2x_x1_3018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv13105_3022,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3041_inst
    process(sext108_3038) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext108_3038(31 downto 0);
      type_cast_3041_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3046_inst
    process(ASHR_i32_i32_3045_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3045_wire(31 downto 0);
      shr_3047 <= tmp_var; -- 
    end process;
    type_cast_3051_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3051_inst_req_0;
      type_cast_3051_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3051_inst_req_1;
      type_cast_3051_inst_ack_1<= rack(0);
      type_cast_3051_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3051_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3050_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom_3052,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_3072_inst
    process(sext109_3069) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := sext109_3069(31 downto 0);
      type_cast_3072_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_3077_inst
    process(ASHR_i32_i32_3076_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := ASHR_i32_i32_3076_wire(31 downto 0);
      shr64_3078 <= tmp_var; -- 
    end process;
    type_cast_3082_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3082_inst_req_0;
      type_cast_3082_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3082_inst_req_1;
      type_cast_3082_inst_ack_1<= rack(0);
      type_cast_3082_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3082_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3081_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => idxprom65_3083,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3098_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3098_inst_req_0;
      type_cast_3098_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3098_inst_req_1;
      type_cast_3098_inst_ack_1<= rack(0);
      type_cast_3098_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3098_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3097_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv69_3099,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3135_inst_req_0;
      type_cast_3135_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3135_inst_req_1;
      type_cast_3135_inst_ack_1<= rack(0);
      type_cast_3135_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3134_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_3136,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3163_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3163_inst_req_0;
      type_cast_3163_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3163_inst_req_1;
      type_cast_3163_inst_ack_1<= rack(0);
      type_cast_3163_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3163_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => div87_3160,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv88_3164,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3170_inst_req_0;
      type_cast_3170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3170_inst_req_1;
      type_cast_3170_inst_ack_1<= rack(0);
      type_cast_3170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv88_3164,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3170_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3172_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3172_inst_req_0;
      type_cast_3172_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3172_inst_req_1;
      type_cast_3172_inst_ack_1<= rack(0);
      type_cast_3172_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3172_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc_3131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3172_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3176_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3176_inst_req_0;
      type_cast_3176_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3176_inst_req_1;
      type_cast_3176_inst_ack_1<= rack(0);
      type_cast_3176_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3176_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inc85_3154,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3176_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3178_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3178_inst_req_0;
      type_cast_3178_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3178_inst_req_1;
      type_cast_3178_inst_ack_1<= rack(0);
      type_cast_3178_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3178_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => input_dim0x_x2x_xph_2884,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_3178_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_3183_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_3183_inst_req_0;
      type_cast_3183_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_3183_inst_req_1;
      type_cast_3183_inst_ack_1<= rack(0);
      type_cast_3183_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_3183_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => type_cast_3182_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv90_3184,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence LOAD_padding_2820_gather_scatter
    process(LOAD_padding_2820_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := LOAD_padding_2820_data_0;
      ov(15 downto 0) := iv;
      tmp30_2821 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3057_index_1_rename
    process(R_idxprom_3056_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom_3056_resized;
      ov(13 downto 0) := iv;
      R_idxprom_3056_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3057_index_1_resize
    process(idxprom_3052) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom_3052;
      ov := iv(13 downto 0);
      R_idxprom_3056_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3057_root_address_inst
    process(array_obj_ref_3057_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3057_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3057_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3088_index_1_rename
    process(R_idxprom65_3087_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_idxprom65_3087_resized;
      ov(13 downto 0) := iv;
      R_idxprom65_3087_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3088_index_1_resize
    process(idxprom65_3083) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := idxprom65_3083;
      ov := iv(13 downto 0);
      R_idxprom65_3087_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_3088_root_address_inst
    process(array_obj_ref_3088_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_3088_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_3088_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2747_addr_0
    process(ptr_deref_2747_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2747_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2747_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2747_base_resize
    process(iNsTr_2_2744) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_2744;
      ov := iv(6 downto 0);
      ptr_deref_2747_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2747_gather_scatter
    process(ptr_deref_2747_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2747_data_0;
      ov(31 downto 0) := iv;
      tmp_2748 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2747_root_address_inst
    process(ptr_deref_2747_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2747_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2747_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2769_addr_0
    process(ptr_deref_2769_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2769_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2769_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2769_base_resize
    process(iNsTr_3_2766) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_3_2766;
      ov := iv(6 downto 0);
      ptr_deref_2769_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2769_gather_scatter
    process(ptr_deref_2769_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2769_data_0;
      ov(31 downto 0) := iv;
      tmp2_2770 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2769_root_address_inst
    process(ptr_deref_2769_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2769_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2769_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_addr_0
    process(ptr_deref_2791_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2791_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_base_resize
    process(iNsTr_4_2788) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_4_2788;
      ov := iv(6 downto 0);
      ptr_deref_2791_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_gather_scatter
    process(ptr_deref_2791_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_data_0;
      ov(31 downto 0) := iv;
      tmp14_2792 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2791_root_address_inst
    process(ptr_deref_2791_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2791_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2791_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2801_addr_0
    process(ptr_deref_2801_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2801_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2801_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2801_base_resize
    process(iNsTr_5_2798) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_2798;
      ov := iv(0 downto 0);
      ptr_deref_2801_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2801_gather_scatter
    process(ptr_deref_2801_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2801_data_0;
      ov(15 downto 0) := iv;
      tmp25_2802 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2801_root_address_inst
    process(ptr_deref_2801_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2801_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2801_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_addr_0
    process(ptr_deref_2817_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2817_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_base_resize
    process(iNsTr_6_2814) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_6_2814;
      ov := iv(6 downto 0);
      ptr_deref_2817_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_gather_scatter
    process(ptr_deref_2817_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_data_0;
      ov(31 downto 0) := iv;
      tmp28_2818 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2817_root_address_inst
    process(ptr_deref_2817_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2817_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2817_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_addr_0
    process(ptr_deref_2834_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2834_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_2834_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_base_resize
    process(iNsTr_7_2831) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_7_2831;
      ov := iv(0 downto 0);
      ptr_deref_2834_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_gather_scatter
    process(ptr_deref_2834_data_0) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2834_data_0;
      ov(15 downto 0) := iv;
      tmp36_2835 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2834_root_address_inst
    process(ptr_deref_2834_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2834_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_2834_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2850_addr_0
    process(ptr_deref_2850_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2850_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2850_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2850_base_resize
    process(iNsTr_8_2847) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_8_2847;
      ov := iv(6 downto 0);
      ptr_deref_2850_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2850_gather_scatter
    process(ptr_deref_2850_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2850_data_0;
      ov(31 downto 0) := iv;
      tmp39_2851 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2850_root_address_inst
    process(ptr_deref_2850_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2850_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2850_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2862_addr_0
    process(ptr_deref_2862_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2862_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2862_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2862_base_resize
    process(iNsTr_9_2859) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_9_2859;
      ov := iv(6 downto 0);
      ptr_deref_2862_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2862_gather_scatter
    process(ptr_deref_2862_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2862_data_0;
      ov(31 downto 0) := iv;
      tmp48_2863 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2862_root_address_inst
    process(ptr_deref_2862_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2862_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2862_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2874_addr_0
    process(ptr_deref_2874_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2874_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_2874_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2874_base_resize
    process(iNsTr_10_2871) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_10_2871;
      ov := iv(6 downto 0);
      ptr_deref_2874_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2874_gather_scatter
    process(ptr_deref_2874_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2874_data_0;
      ov(31 downto 0) := iv;
      tmp51_2875 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_2874_root_address_inst
    process(ptr_deref_2874_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_2874_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_2874_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3062_addr_0
    process(ptr_deref_3062_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3062_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3062_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3062_base_resize
    process(arrayidx_3059) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_3059;
      ov := iv(13 downto 0);
      ptr_deref_3062_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3062_gather_scatter
    process(ptr_deref_3062_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3062_data_0;
      ov(63 downto 0) := iv;
      tmp61_3063 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3062_root_address_inst
    process(ptr_deref_3062_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3062_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3062_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_addr_0
    process(ptr_deref_3092_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3092_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_3092_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_base_resize
    process(arrayidx66_3090) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx66_3090;
      ov := iv(13 downto 0);
      ptr_deref_3092_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_gather_scatter
    process(tmp61_3063) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := tmp61_3063;
      ov(63 downto 0) := iv;
      ptr_deref_3092_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_3092_root_address_inst
    process(ptr_deref_3092_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_3092_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_3092_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_3111_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_3110;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3111_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3111_branch_req_0,
          ack0 => if_stmt_3111_branch_ack_0,
          ack1 => if_stmt_3111_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3142_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp81_3141;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3142_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3142_branch_req_0,
          ack0 => if_stmt_3142_branch_ack_0,
          ack1 => if_stmt_3142_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3190_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp92_3189;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3190_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3190_branch_req_0,
          ack0 => if_stmt_3190_branch_ack_0,
          ack1 => if_stmt_3190_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u16_u16_3122_inst
    process(indvar_3005) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_3005, type_cast_3121_wire_constant, tmp_var);
      indvarx_xnext_3123 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3130_inst
    process(input_dim1x_x1x_xph_2878) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim1x_x1x_xph_2878, type_cast_3129_wire_constant, tmp_var);
      inc_3131 <= tmp_var; --
    end process;
    -- binary operator ADD_u16_u16_3153_inst
    process(input_dim0x_x2x_xph_2884) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntAdd_proc(input_dim0x_x2x_xph_2884, type_cast_3152_wire_constant, tmp_var);
      inc85_3154 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2909_inst
    process(mul_2905, conv16_2895) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul_2905, conv16_2895, tmp_var);
      add_2910 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2924_inst
    process(mul27_2920, tmp28_2818) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul27_2920, tmp28_2818, tmp_var);
      add29_2925 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2939_inst
    process(mul38_2935, tmp39_2851) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul38_2935, tmp39_2851, tmp_var);
      add40_2940 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2956_inst
    process(sub44_2951) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub44_2951, type_cast_2955_wire_constant, tmp_var);
      sext_2957 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2977_inst
    process(sub32_2972) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(sub32_2972, type_cast_2976_wire_constant, tmp_var);
      sext106_2978 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_2996_inst
    process(conv50_2966, mul54_2992) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv50_2966, mul54_2992, tmp_var);
      add55_2997 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3026_inst
    process(mul20_2915, conv13105_3022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul20_2915, conv13105_3022, tmp_var);
      add21_3027 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3031_inst
    process(mul56_3002, conv13105_3022) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mul56_3002, conv13105_3022, tmp_var);
      add57_3032 <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_3104_inst
    process(conv69_3099) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(conv69_3099, type_cast_3103_wire_constant, tmp_var);
      add70_3105 <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2964_inst
    process(type_cast_2960_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2960_wire, type_cast_2963_wire_constant, tmp_var);
      ASHR_i32_i32_2964_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_2985_inst
    process(type_cast_2981_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_2981_wire, type_cast_2984_wire_constant, tmp_var);
      ASHR_i32_i32_2985_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3045_inst
    process(type_cast_3041_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3041_wire, type_cast_3044_wire_constant, tmp_var);
      ASHR_i32_i32_3045_wire <= tmp_var; --
    end process;
    -- binary operator ASHR_i32_i32_3076_inst
    process(type_cast_3072_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntASHR_proc(type_cast_3072_wire, type_cast_3075_wire_constant, tmp_var);
      ASHR_i32_i32_3076_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3140_inst
    process(conv79_3136, tmp2_2770) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv79_3136, tmp2_2770, tmp_var);
      cmp81_3141 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_3188_inst
    process(conv90_3184, tmp_2748) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv90_3184, tmp_2748, tmp_var);
      cmp92_3189 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2753_inst
    process(tmp_2748) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp_2748, type_cast_2752_wire_constant, tmp_var);
      div_2754 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_2775_inst
    process(tmp2_2770) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2770, type_cast_2774_wire_constant, tmp_var);
      div3_2776 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_3159_inst
    process(tmp2_2770) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp2_2770, type_cast_3158_wire_constant, tmp_var);
      div87_3160 <= tmp_var; --
    end process;
    -- binary operator MUL_u16_u16_3017_inst
    process(indvar_3005) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntMul_proc(indvar_3005, type_cast_3016_wire_constant, tmp_var);
      input_dim2x_x1_3018 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2904_inst
    process(tmp2_2770, conv19_2900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp2_2770, conv19_2900, tmp_var);
      mul_2905 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2914_inst
    process(add_2910, tmp14_2792) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add_2910, tmp14_2792, tmp_var);
      mul20_2915 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2919_inst
    process(conv26_2806, conv19_2900) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv26_2806, conv19_2900, tmp_var);
      mul27_2920 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2934_inst
    process(conv37_2839, conv16_2895) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(conv37_2839, conv16_2895, tmp_var);
      mul38_2935 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_2991_inst
    process(tmp51_2875, conv53_2987) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp51_2875, conv53_2987, tmp_var);
      mul54_2992 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_3001_inst
    process(add55_2997, tmp48_2863) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(add55_2997, tmp48_2863, tmp_var);
      mul56_3002 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2950_inst
    process(sub43_2945) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub43_2945, type_cast_2949_wire_constant, tmp_var);
      sub44_2951 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_2971_inst
    process(sub_2930) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(sub_2930, type_cast_2970_wire_constant, tmp_var);
      sub32_2972 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3037_inst
    process(add21_3027) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add21_3027, type_cast_3036_wire_constant, tmp_var);
      sext108_3038 <= tmp_var; --
    end process;
    -- binary operator SHL_u32_u32_3068_inst
    process(add57_3032) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add57_3032, type_cast_3067_wire_constant, tmp_var);
      sext109_3069 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2929_inst
    process(add29_2925, conv31_2825) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add29_2925, conv31_2825, tmp_var);
      sub_2930 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_2944_inst
    process(add40_2940, conv31_2825) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(add40_2940, conv31_2825, tmp_var);
      sub43_2945 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_3109_inst
    process(add70_3105, tmp14_2792) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(add70_3105, tmp14_2792, tmp_var);
      cmp_3110 <= tmp_var; --
    end process;
    -- shared split operator group (35) : array_obj_ref_3057_index_offset 
    ApIntAdd_group_35: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom_3056_scaled;
      array_obj_ref_3057_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3057_index_offset_req_0;
      array_obj_ref_3057_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3057_index_offset_req_1;
      array_obj_ref_3057_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_35_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_35_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_35",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : array_obj_ref_3088_index_offset 
    ApIntAdd_group_36: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_idxprom65_3087_scaled;
      array_obj_ref_3088_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_3088_index_offset_req_0;
      array_obj_ref_3088_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_3088_index_offset_req_1;
      array_obj_ref_3088_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_36_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_36_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_36",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- unary operator type_cast_2893_inst
    process(input_dim1x_x1x_xph_2878) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim1x_x1x_xph_2878, tmp_var);
      type_cast_2893_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_2898_inst
    process(input_dim0x_x2x_xph_2884) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x2x_xph_2884, tmp_var);
      type_cast_2898_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3050_inst
    process(shr_3047) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr_3047, tmp_var);
      type_cast_3050_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3081_inst
    process(shr64_3078) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", shr64_3078, tmp_var);
      type_cast_3081_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3097_inst
    process(input_dim2x_x1_3018) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim2x_x1_3018, tmp_var);
      type_cast_3097_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3134_inst
    process(inc_3131) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", inc_3131, tmp_var);
      type_cast_3134_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_3182_inst
    process(input_dim0x_x0_3173) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", input_dim0x_x0_3173, tmp_var);
      type_cast_3182_wire <= tmp_var; -- 
    end process;
    -- shared load operator group (0) : LOAD_padding_2820_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= LOAD_padding_2820_load_0_req_0;
      LOAD_padding_2820_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= LOAD_padding_2820_load_0_req_1;
      LOAD_padding_2820_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= LOAD_padding_2820_word_address_0;
      LOAD_padding_2820_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(15 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_2747_load_0 ptr_deref_2769_load_0 ptr_deref_2791_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_2747_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_2769_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2791_load_0_req_0;
      ptr_deref_2747_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_2769_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2791_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_2747_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_2769_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2791_load_0_req_1;
      ptr_deref_2747_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_2769_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2791_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2747_word_address_0 & ptr_deref_2769_word_address_0 & ptr_deref_2791_word_address_0;
      ptr_deref_2747_data_0 <= data_out(95 downto 64);
      ptr_deref_2769_data_0 <= data_out(63 downto 32);
      ptr_deref_2791_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 3,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2801_load_0 ptr_deref_2834_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2801_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2834_load_0_req_0;
      ptr_deref_2801_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2834_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2801_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2834_load_0_req_1;
      ptr_deref_2801_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2834_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2801_word_address_0 & ptr_deref_2834_word_address_0;
      ptr_deref_2801_data_0 <= data_out(31 downto 16);
      ptr_deref_2834_data_0 <= data_out(15 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 16,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(15 downto 0),
          mtag => memory_space_7_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2817_load_0 ptr_deref_2850_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2817_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2850_load_0_req_0;
      ptr_deref_2817_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2850_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2817_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2850_load_0_req_1;
      ptr_deref_2817_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2850_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup3_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup3_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup3_gI: SplitGuardInterface generic map(name => "LoadGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2817_word_address_0 & ptr_deref_2850_word_address_0;
      ptr_deref_2817_data_0 <= data_out(63 downto 32);
      ptr_deref_2850_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup3", addr_width => 7,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup3 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2862_load_0 ptr_deref_2874_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_2862_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_2874_load_0_req_0;
      ptr_deref_2862_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_2874_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_2862_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_2874_load_0_req_1;
      ptr_deref_2862_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_2874_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      LoadGroup4_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup4_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup4_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup4_gI: SplitGuardInterface generic map(name => "LoadGroup4_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_2862_word_address_0 & ptr_deref_2874_word_address_0;
      ptr_deref_2862_data_0 <= data_out(63 downto 32);
      ptr_deref_2874_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup4", addr_width => 7,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup4 load-complete ",
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_3062_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3062_load_0_req_0;
      ptr_deref_3062_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3062_load_0_req_1;
      ptr_deref_3062_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup5_gI: SplitGuardInterface generic map(name => "LoadGroup5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_3062_word_address_0;
      ptr_deref_3062_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup5", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup5 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(63 downto 0),
          mtag => memory_space_3_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared store operator group (0) : ptr_deref_3092_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_3092_store_0_req_0;
      ptr_deref_3092_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_3092_store_0_req_1;
      ptr_deref_3092_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_3092_word_address_0;
      data_in <= ptr_deref_3092_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_Block3_start_2734_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_Block3_start_2734_inst_req_0;
      RPIPE_Block3_start_2734_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_Block3_start_2734_inst_req_1;
      RPIPE_Block3_start_2734_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      call_2735 <= data_out(15 downto 0);
      Block3_start_read_0_gI: SplitGuardInterface generic map(name => "Block3_start_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      Block3_start_read_0: InputPortRevised -- 
        generic map ( name => "Block3_start_read_0", data_width => 16,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => Block3_start_pipe_read_req(0),
          oack => Block3_start_pipe_read_ack(0),
          odata => Block3_start_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_Block3_done_3198_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_Block3_done_3198_inst_req_0;
      WPIPE_Block3_done_3198_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_Block3_done_3198_inst_req_1;
      WPIPE_Block3_done_3198_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= call_2735;
      Block3_done_write_0_gI: SplitGuardInterface generic map(name => "Block3_done_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      Block3_done_write_0: OutputPortRevised -- 
        generic map ( name => "Block3_done", data_width => 16, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => Block3_done_pipe_write_req(0),
          oack => Block3_done_pipe_write_ack(0),
          odata => Block3_done_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end convTransposeD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity sendOutput is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sendOutput;
architecture sendOutput_arch of sendOutput is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal sendOutput_CP_3266_start: Boolean;
  signal sendOutput_CP_3266_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal array_obj_ref_1199_index_offset_ack_0 : boolean;
  signal ptr_deref_1113_load_0_req_1 : boolean;
  signal ptr_deref_1113_load_0_ack_0 : boolean;
  signal type_cast_1170_inst_ack_0 : boolean;
  signal ptr_deref_1113_load_0_ack_1 : boolean;
  signal type_cast_1170_inst_req_0 : boolean;
  signal array_obj_ref_1199_index_offset_req_1 : boolean;
  signal array_obj_ref_1199_index_offset_ack_1 : boolean;
  signal array_obj_ref_1199_index_offset_req_0 : boolean;
  signal ptr_deref_1113_load_0_req_0 : boolean;
  signal ptr_deref_1101_load_0_ack_1 : boolean;
  signal addr_of_1200_final_reg_req_1 : boolean;
  signal ptr_deref_1101_load_0_req_1 : boolean;
  signal type_cast_1208_inst_ack_0 : boolean;
  signal type_cast_1228_inst_req_0 : boolean;
  signal ptr_deref_1101_load_0_ack_0 : boolean;
  signal type_cast_1228_inst_req_1 : boolean;
  signal type_cast_1218_inst_ack_1 : boolean;
  signal type_cast_1238_inst_req_0 : boolean;
  signal type_cast_1238_inst_req_1 : boolean;
  signal type_cast_1170_inst_req_1 : boolean;
  signal type_cast_1218_inst_req_1 : boolean;
  signal type_cast_1258_inst_req_1 : boolean;
  signal type_cast_1170_inst_ack_1 : boolean;
  signal ptr_deref_1204_load_0_req_0 : boolean;
  signal ptr_deref_1125_load_0_req_1 : boolean;
  signal type_cast_1208_inst_req_1 : boolean;
  signal type_cast_1268_inst_req_1 : boolean;
  signal type_cast_1268_inst_ack_1 : boolean;
  signal type_cast_1208_inst_ack_1 : boolean;
  signal addr_of_1200_final_reg_req_0 : boolean;
  signal type_cast_1228_inst_ack_1 : boolean;
  signal type_cast_1238_inst_ack_0 : boolean;
  signal ptr_deref_1204_load_0_ack_0 : boolean;
  signal addr_of_1200_final_reg_ack_0 : boolean;
  signal type_cast_1268_inst_req_0 : boolean;
  signal type_cast_1268_inst_ack_0 : boolean;
  signal type_cast_1228_inst_ack_0 : boolean;
  signal type_cast_1248_inst_req_1 : boolean;
  signal addr_of_1200_final_reg_ack_1 : boolean;
  signal ptr_deref_1101_load_0_req_0 : boolean;
  signal type_cast_1248_inst_req_0 : boolean;
  signal type_cast_1258_inst_ack_1 : boolean;
  signal ptr_deref_1125_load_0_req_0 : boolean;
  signal ptr_deref_1125_load_0_ack_0 : boolean;
  signal ptr_deref_1125_load_0_ack_1 : boolean;
  signal type_cast_1238_inst_ack_1 : boolean;
  signal type_cast_1218_inst_req_0 : boolean;
  signal type_cast_1208_inst_req_0 : boolean;
  signal type_cast_1248_inst_ack_1 : boolean;
  signal ptr_deref_1204_load_0_ack_1 : boolean;
  signal if_stmt_1143_branch_ack_0 : boolean;
  signal if_stmt_1143_branch_ack_1 : boolean;
  signal if_stmt_1143_branch_req_0 : boolean;
  signal type_cast_1218_inst_ack_0 : boolean;
  signal ptr_deref_1204_load_0_req_1 : boolean;
  signal type_cast_1248_inst_ack_0 : boolean;
  signal type_cast_1258_inst_req_0 : boolean;
  signal type_cast_1258_inst_ack_0 : boolean;
  signal type_cast_1278_inst_req_0 : boolean;
  signal type_cast_1278_inst_ack_0 : boolean;
  signal type_cast_1278_inst_req_1 : boolean;
  signal type_cast_1278_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_req_1 : boolean;
  signal WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 : boolean;
  signal if_stmt_1315_branch_req_0 : boolean;
  signal if_stmt_1315_branch_ack_1 : boolean;
  signal if_stmt_1315_branch_ack_0 : boolean;
  signal phi_stmt_1187_req_0 : boolean;
  signal type_cast_1193_inst_req_0 : boolean;
  signal type_cast_1193_inst_ack_0 : boolean;
  signal type_cast_1193_inst_req_1 : boolean;
  signal type_cast_1193_inst_ack_1 : boolean;
  signal phi_stmt_1187_req_1 : boolean;
  signal phi_stmt_1187_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "sendOutput_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  sendOutput_CP_3266_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "sendOutput_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3266_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sendOutput_CP_3266_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= sendOutput_CP_3266_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  sendOutput_CP_3266: Block -- control-path 
    signal sendOutput_CP_3266_elements: BooleanArray(66 downto 0);
    -- 
  begin -- 
    sendOutput_CP_3266_elements(0) <= sendOutput_CP_3266_start;
    sendOutput_CP_3266_symbol <= sendOutput_CP_3266_elements(66);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	6 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (83) 
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142__entry__
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/branch_block_stmt_1090__entry__
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/word_0/rr
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/$entry
      -- CP-element group 0: 	 branch_block_stmt_1090/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_update_start_
      -- CP-element group 0: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_base_addr_resize/$entry
      -- 
    cr_3390_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3390_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1113_load_0_req_1); -- 
    rr_3379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1113_load_0_req_0); -- 
    cr_3340_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3340_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1101_load_0_req_1); -- 
    cr_3440_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3440_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1125_load_0_req_1); -- 
    rr_3329_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3329_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1101_load_0_req_0); -- 
    rr_3429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(0), ack => ptr_deref_1125_load_0_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/word_0/ra
      -- CP-element group 1: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_sample_completed_
      -- 
    ra_3330_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1101_load_0_ack_0, ack => sendOutput_CP_3266_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/ptr_deref_1101_Merge/$entry
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/ptr_deref_1101_Merge/merge_ack
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/ptr_deref_1101_Merge/merge_req
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/ptr_deref_1101_Merge/$exit
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1101_update_completed_
      -- 
    ca_3341_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1101_load_0_ack_1, ack => sendOutput_CP_3266_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (5) 
      -- CP-element group 3: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/word_0/ra
      -- CP-element group 3: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/word_0/$exit
      -- CP-element group 3: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/word_access_start/$exit
      -- CP-element group 3: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Sample/$exit
      -- 
    ra_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_0, ack => sendOutput_CP_3266_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (9) 
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/ptr_deref_1113_Merge/$exit
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/word_0/$exit
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/word_access_complete/word_0/ca
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/ptr_deref_1113_Merge/$entry
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/ptr_deref_1113_Merge/merge_req
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_Update/ptr_deref_1113_Merge/merge_ack
      -- CP-element group 4: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1113_update_completed_
      -- 
    ca_3391_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1113_load_0_ack_1, ack => sendOutput_CP_3266_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/$exit
      -- CP-element group 5: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/word_0/$exit
      -- CP-element group 5: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Sample/word_access_start/word_0/ra
      -- CP-element group 5: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_sample_completed_
      -- 
    ra_3430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_0, ack => sendOutput_CP_3266_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	0 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (9) 
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/$exit
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/ptr_deref_1125_Merge/merge_req
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/ptr_deref_1125_Merge/merge_ack
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/word_access_complete/word_0/ca
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/ptr_deref_1125_Merge/$exit
      -- CP-element group 6: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/ptr_deref_1125_Update/ptr_deref_1125_Merge/$entry
      -- 
    ca_3441_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1125_load_0_ack_1, ack => sendOutput_CP_3266_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (10) 
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143__entry__
      -- CP-element group 7: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142__exit__
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_eval_test/$exit
      -- CP-element group 7: 	 branch_block_stmt_1090/assign_stmt_1098_to_assign_stmt_1142/$exit
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_else_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_1090/R_cmp73_1144_place
      -- CP-element group 7: 	 branch_block_stmt_1090/if_stmt_1143_eval_test/branch_req
      -- 
    branch_req_3454_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3454_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(7), ack => if_stmt_1143_branch_req_0); -- 
    sendOutput_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "sendOutput_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(4) & sendOutput_CP_3266_elements(2) & sendOutput_CP_3266_elements(6);
      gj_sendOutput_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (18) 
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_update_start_
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184__entry__
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Sample/rr
      -- CP-element group 8: 	 branch_block_stmt_1090/merge_stmt_1149__exit__
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_sample_start_
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Update/cr
      -- CP-element group 8: 	 branch_block_stmt_1090/entry_bbx_xnph
      -- CP-element group 8: 	 branch_block_stmt_1090/if_stmt_1143_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_1090/if_stmt_1143_if_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/$entry
      -- CP-element group 8: 	 branch_block_stmt_1090/entry_bbx_xnph_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_1090/entry_bbx_xnph_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_1090/merge_stmt_1149_PhiReqMerge
      -- CP-element group 8: 	 branch_block_stmt_1090/merge_stmt_1149_PhiAck/$entry
      -- CP-element group 8: 	 branch_block_stmt_1090/merge_stmt_1149_PhiAck/$exit
      -- CP-element group 8: 	 branch_block_stmt_1090/merge_stmt_1149_PhiAck/dummy
      -- 
    if_choice_transition_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1143_branch_ack_1, ack => sendOutput_CP_3266_elements(8)); -- 
    rr_3476_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3476_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(8), ack => type_cast_1170_inst_req_0); -- 
    cr_3481_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3481_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(8), ack => type_cast_1170_inst_req_1); -- 
    -- CP-element group 9:  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	66 
    -- CP-element group 9:  members (5) 
      -- CP-element group 9: 	 branch_block_stmt_1090/entry_forx_xend
      -- CP-element group 9: 	 branch_block_stmt_1090/if_stmt_1143_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_1090/if_stmt_1143_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_1090/entry_forx_xend_PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_1090/entry_forx_xend_PhiReq/$exit
      -- 
    else_choice_transition_3463_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1143_branch_ack_0, ack => sendOutput_CP_3266_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Sample/ra
      -- CP-element group 10: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_sample_completed_
      -- 
    ra_3477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1170_inst_ack_0, ack => sendOutput_CP_3266_elements(10)); -- 
    -- CP-element group 11:  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	60 
    -- CP-element group 11:  members (9) 
      -- CP-element group 11: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody
      -- CP-element group 11: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184__exit__
      -- CP-element group 11: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/type_cast_1170_Update/ca
      -- CP-element group 11: 	 branch_block_stmt_1090/assign_stmt_1155_to_assign_stmt_1184/$exit
      -- CP-element group 11: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/$entry
      -- CP-element group 11: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/$entry
      -- CP-element group 11: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/$entry
      -- 
    ca_3482_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1170_inst_ack_1, ack => sendOutput_CP_3266_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	65 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	57 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Sample/ack
      -- CP-element group 12: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_sample_complete
      -- 
    ack_3511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1199_index_offset_ack_0, ack => sendOutput_CP_3266_elements(12)); -- 
    -- CP-element group 13:  transition  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	65 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (11) 
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_base_plus_offset/$exit
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_root_address_calculated
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_base_plus_offset/$entry
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Update/ack
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_base_plus_offset/sum_rename_req
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_base_plus_offset/sum_rename_ack
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_request/$entry
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_offset_calculated
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_request/req
      -- CP-element group 13: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_sample_start_
      -- 
    ack_3516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1199_index_offset_ack_1, ack => sendOutput_CP_3266_elements(13)); -- 
    req_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(13), ack => addr_of_1200_final_reg_req_0); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_request/$exit
      -- CP-element group 14: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_request/ack
      -- CP-element group 14: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_sample_completed_
      -- 
    ack_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1200_final_reg_ack_0, ack => sendOutput_CP_3266_elements(14)); -- 
    -- CP-element group 15:  join  fork  transition  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	65 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (24) 
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_complete/$exit
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_address_resized
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_addr_resize/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_addr_resize/$exit
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_complete/ack
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_addr_resize/base_resize_req
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_base_addr_resize/base_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_word_address_calculated
      -- 
    ack_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1200_final_reg_ack_1, ack => sendOutput_CP_3266_elements(15)); -- 
    rr_3564_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3564_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(15), ack => ptr_deref_1204_load_0_req_0); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (5) 
      -- CP-element group 16: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/$exit
      -- CP-element group 16: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/word_0/$exit
      -- CP-element group 16: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Sample/word_access_start/word_0/ra
      -- 
    ra_3565_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1204_load_0_ack_0, ack => sendOutput_CP_3266_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	65 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	32 
    -- CP-element group 17: 	18 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	28 
    -- CP-element group 17: 	30 
    -- CP-element group 17: 	26 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	22 
    -- CP-element group 17:  members (33) 
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/ptr_deref_1204_Merge/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/ptr_deref_1204_Merge/$exit
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/$exit
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/ptr_deref_1204_Merge/merge_req
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/ptr_deref_1204_Merge/merge_ack
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/word_0/$exit
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_sample_start_
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/word_0/ca
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Sample/rr
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Sample/$entry
      -- CP-element group 17: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Sample/rr
      -- 
    ca_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1204_load_0_ack_1, ack => sendOutput_CP_3266_elements(17)); -- 
    rr_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1278_inst_req_0); -- 
    rr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1218_inst_req_0); -- 
    rr_3589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1208_inst_req_0); -- 
    rr_3673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1268_inst_req_0); -- 
    rr_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1258_inst_req_0); -- 
    rr_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1238_inst_req_0); -- 
    rr_3645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1248_inst_req_0); -- 
    rr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(17), ack => type_cast_1228_inst_req_0); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_sample_completed_
      -- CP-element group 18: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Sample/ra
      -- CP-element group 18: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Sample/$exit
      -- 
    ra_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_0, ack => sendOutput_CP_3266_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	65 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	54 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Update/ca
      -- 
    ca_3595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1208_inst_ack_1, ack => sendOutput_CP_3266_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	17 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_sample_completed_
      -- CP-element group 20: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Sample/ra
      -- CP-element group 20: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Sample/$exit
      -- 
    ra_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_0, ack => sendOutput_CP_3266_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	65 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	51 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Update/ca
      -- CP-element group 21: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_update_completed_
      -- CP-element group 21: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Update/$exit
      -- 
    ca_3609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1218_inst_ack_1, ack => sendOutput_CP_3266_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	17 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Sample/ra
      -- CP-element group 22: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Sample/$exit
      -- 
    ra_3618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_0, ack => sendOutput_CP_3266_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	48 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Update/ca
      -- 
    ca_3623_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1228_inst_ack_1, ack => sendOutput_CP_3266_elements(23)); -- 
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	17 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Sample/ra
      -- 
    ra_3632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_0, ack => sendOutput_CP_3266_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	65 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	45 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Update/ca
      -- 
    ca_3637_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1238_inst_ack_1, ack => sendOutput_CP_3266_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	17 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Sample/ra
      -- 
    ra_3646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_0, ack => sendOutput_CP_3266_elements(26)); -- 
    -- CP-element group 27:  transition  input  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	65 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	42 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_update_completed_
      -- 
    ca_3651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1248_inst_ack_1, ack => sendOutput_CP_3266_elements(27)); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	17 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Sample/ra
      -- CP-element group 28: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Sample/$exit
      -- 
    ra_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_0, ack => sendOutput_CP_3266_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	65 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	39 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Update/ca
      -- CP-element group 29: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_update_completed_
      -- 
    ca_3665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1258_inst_ack_1, ack => sendOutput_CP_3266_elements(29)); -- 
    -- CP-element group 30:  transition  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	17 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_sample_completed_
      -- 
    ra_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1268_inst_ack_0, ack => sendOutput_CP_3266_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	65 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	36 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_update_completed_
      -- CP-element group 31: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Update/ca
      -- 
    ca_3679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1268_inst_ack_1, ack => sendOutput_CP_3266_elements(31)); -- 
    -- CP-element group 32:  transition  input  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	17 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Sample/ra
      -- 
    ra_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1278_inst_ack_0, ack => sendOutput_CP_3266_elements(32)); -- 
    -- CP-element group 33:  transition  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	65 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	34 
    -- CP-element group 33:  members (6) 
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Update/ca
      -- CP-element group 33: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Sample/req
      -- 
    ca_3693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1278_inst_ack_1, ack => sendOutput_CP_3266_elements(33)); -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(33), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_0); -- 
    -- CP-element group 34:  transition  input  output  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	33 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	35 
    -- CP-element group 34:  members (6) 
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_update_start_
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Update/req
      -- 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0, ack => sendOutput_CP_3266_elements(34)); -- 
    req_3706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(34), ack => WPIPE_ConvTranspose_output_pipe_1280_inst_req_1); -- 
    -- CP-element group 35:  transition  input  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	34 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1280_Update/ack
      -- 
    ack_3707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1, ack => sendOutput_CP_3266_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: 	31 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	37 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_sample_start_
      -- CP-element group 36: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Sample/req
      -- 
    req_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(36), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_0); -- 
    sendOutput_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(35) & sendOutput_CP_3266_elements(31);
      gj_sendOutput_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  transition  input  output  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	38 
    -- CP-element group 37:  members (6) 
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_update_start_
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Sample/ack
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Update/$entry
      -- CP-element group 37: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Update/req
      -- 
    ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0, ack => sendOutput_CP_3266_elements(37)); -- 
    req_3720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(37), ack => WPIPE_ConvTranspose_output_pipe_1283_inst_req_1); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	39 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1283_Update/ack
      -- 
    ack_3721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1, ack => sendOutput_CP_3266_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	29 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Sample/req
      -- 
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(39), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_0); -- 
    sendOutput_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(38) & sendOutput_CP_3266_elements(29);
      gj_sendOutput_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  transition  input  output  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	39 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	41 
    -- CP-element group 40:  members (6) 
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Sample/ack
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Update/req
      -- 
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0, ack => sendOutput_CP_3266_elements(40)); -- 
    req_3734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(40), ack => WPIPE_ConvTranspose_output_pipe_1286_inst_req_1); -- 
    -- CP-element group 41:  transition  input  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	40 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1286_Update/ack
      -- 
    ack_3735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1, ack => sendOutput_CP_3266_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	27 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	43 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Sample/req
      -- 
    req_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(42), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_0); -- 
    sendOutput_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(41) & sendOutput_CP_3266_elements(27);
      gj_sendOutput_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  transition  input  output  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	42 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	44 
    -- CP-element group 43:  members (6) 
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Sample/ack
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Update/req
      -- 
    ack_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0, ack => sendOutput_CP_3266_elements(43)); -- 
    req_3748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(43), ack => WPIPE_ConvTranspose_output_pipe_1289_inst_req_1); -- 
    -- CP-element group 44:  transition  input  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	43 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1289_Update/ack
      -- 
    ack_3749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1, ack => sendOutput_CP_3266_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: 	25 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Sample/req
      -- 
    req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(45), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_0); -- 
    sendOutput_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(44) & sendOutput_CP_3266_elements(25);
      gj_sendOutput_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  transition  input  output  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	47 
    -- CP-element group 46:  members (6) 
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Update/req
      -- 
    ack_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0, ack => sendOutput_CP_3266_elements(46)); -- 
    req_3762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(46), ack => WPIPE_ConvTranspose_output_pipe_1292_inst_req_1); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	46 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1292_Update/ack
      -- 
    ack_3763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1, ack => sendOutput_CP_3266_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	23 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Sample/req
      -- 
    req_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(48), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_0); -- 
    sendOutput_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(47) & sendOutput_CP_3266_elements(23);
      gj_sendOutput_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  output  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	50 
    -- CP-element group 49:  members (6) 
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_update_start_
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Sample/ack
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Update/$entry
      -- CP-element group 49: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Update/req
      -- 
    ack_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0, ack => sendOutput_CP_3266_elements(49)); -- 
    req_3776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(49), ack => WPIPE_ConvTranspose_output_pipe_1295_inst_req_1); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	49 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	51 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1295_Update/ack
      -- 
    ack_3777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1, ack => sendOutput_CP_3266_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	50 
    -- CP-element group 51: 	21 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Sample/req
      -- 
    req_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(51), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_0); -- 
    sendOutput_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(50) & sendOutput_CP_3266_elements(21);
      gj_sendOutput_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  output  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	53 
    -- CP-element group 52:  members (6) 
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_update_start_
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Sample/ack
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Update/req
      -- 
    ack_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0, ack => sendOutput_CP_3266_elements(52)); -- 
    req_3790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(52), ack => WPIPE_ConvTranspose_output_pipe_1298_inst_req_1); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	52 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	54 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1298_Update/ack
      -- 
    ack_3791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1, ack => sendOutput_CP_3266_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	19 
    -- CP-element group 54: 	53 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	55 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Sample/req
      -- 
    req_3799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(54), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_0); -- 
    sendOutput_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(19) & sendOutput_CP_3266_elements(53);
      gj_sendOutput_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  transition  input  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	54 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (6) 
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Update/req
      -- 
    ack_3800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0, ack => sendOutput_CP_3266_elements(55)); -- 
    req_3804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(55), ack => WPIPE_ConvTranspose_output_pipe_1301_inst_req_1); -- 
    -- CP-element group 56:  transition  input  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/WPIPE_ConvTranspose_output_pipe_1301_Update/ack
      -- 
    ack_3805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1, ack => sendOutput_CP_3266_elements(56)); -- 
    -- CP-element group 57:  branch  join  transition  place  output  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	56 
    -- CP-element group 57: 	12 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (10) 
      -- CP-element group 57: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314__exit__
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315__entry__
      -- CP-element group 57: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/$exit
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_dead_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_eval_test/$entry
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_eval_test/$exit
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_eval_test/branch_req
      -- CP-element group 57: 	 branch_block_stmt_1090/R_exitcond1_1316_place
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_if_link/$entry
      -- CP-element group 57: 	 branch_block_stmt_1090/if_stmt_1315_else_link/$entry
      -- 
    branch_req_3813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(57), ack => if_stmt_1315_branch_req_0); -- 
    sendOutput_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(56) & sendOutput_CP_3266_elements(12);
      gj_sendOutput_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  merge  transition  place  input  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	66 
    -- CP-element group 58:  members (13) 
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xendx_xloopexit_forx_xend
      -- CP-element group 58: 	 branch_block_stmt_1090/merge_stmt_1321__exit__
      -- CP-element group 58: 	 branch_block_stmt_1090/if_stmt_1315_if_link/$exit
      -- CP-element group 58: 	 branch_block_stmt_1090/if_stmt_1315_if_link/if_choice_transition
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 58: 	 branch_block_stmt_1090/merge_stmt_1321_PhiReqMerge
      -- CP-element group 58: 	 branch_block_stmt_1090/merge_stmt_1321_PhiAck/$entry
      -- CP-element group 58: 	 branch_block_stmt_1090/merge_stmt_1321_PhiAck/$exit
      -- CP-element group 58: 	 branch_block_stmt_1090/merge_stmt_1321_PhiAck/dummy
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 58: 	 branch_block_stmt_1090/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- 
    if_choice_transition_3818_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1315_branch_ack_1, ack => sendOutput_CP_3266_elements(58)); -- 
    -- CP-element group 59:  fork  transition  place  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: 	62 
    -- CP-element group 59:  members (12) 
      -- CP-element group 59: 	 branch_block_stmt_1090/if_stmt_1315_else_link/$exit
      -- CP-element group 59: 	 branch_block_stmt_1090/if_stmt_1315_else_link/else_choice_transition
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Sample/rr
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Update/cr
      -- 
    else_choice_transition_3822_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1315_branch_ack_0, ack => sendOutput_CP_3266_elements(59)); -- 
    rr_3866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(59), ack => type_cast_1193_inst_req_0); -- 
    cr_3871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(59), ack => type_cast_1193_inst_req_1); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	11 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	64 
    -- CP-element group 60:  members (5) 
      -- CP-element group 60: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/$exit
      -- CP-element group 60: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/$exit
      -- CP-element group 60: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/$exit
      -- CP-element group 60: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1191_konst_delay_trans
      -- CP-element group 60: 	 branch_block_stmt_1090/bbx_xnph_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_req
      -- 
    phi_stmt_1187_req_3847_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1187_req_3847_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(60), ack => phi_stmt_1187_req_0); -- 
    -- Element group sendOutput_CP_3266_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => sendOutput_CP_3266_elements(11), ack => sendOutput_CP_3266_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  input  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Sample/ra
      -- 
    ra_3867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1193_inst_ack_0, ack => sendOutput_CP_3266_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	63 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/Update/ca
      -- 
    ca_3872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1193_inst_ack_1, ack => sendOutput_CP_3266_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	62 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (6) 
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/$exit
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/$exit
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/$exit
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/$exit
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_sources/type_cast_1193/SplitProtocol/$exit
      -- CP-element group 63: 	 branch_block_stmt_1090/forx_xbody_forx_xbody_PhiReq/phi_stmt_1187/phi_stmt_1187_req
      -- 
    phi_stmt_1187_req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1187_req_3873_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(63), ack => phi_stmt_1187_req_1); -- 
    sendOutput_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "sendOutput_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= sendOutput_CP_3266_elements(61) & sendOutput_CP_3266_elements(62);
      gj_sendOutput_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => sendOutput_CP_3266_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  merge  transition  place  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: 	60 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1090/merge_stmt_1186_PhiReqMerge
      -- CP-element group 64: 	 branch_block_stmt_1090/merge_stmt_1186_PhiAck/$entry
      -- 
    sendOutput_CP_3266_elements(64) <= OrReduce(sendOutput_CP_3266_elements(63) & sendOutput_CP_3266_elements(60));
    -- CP-element group 65:  fork  transition  place  input  output  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	31 
    -- CP-element group 65: 	33 
    -- CP-element group 65: 	19 
    -- CP-element group 65: 	17 
    -- CP-element group 65: 	12 
    -- CP-element group 65: 	29 
    -- CP-element group 65: 	27 
    -- CP-element group 65: 	13 
    -- CP-element group 65: 	15 
    -- CP-element group 65: 	25 
    -- CP-element group 65: 	21 
    -- CP-element group 65: 	23 
    -- CP-element group 65:  members (53) 
      -- CP-element group 65: 	 branch_block_stmt_1090/merge_stmt_1186__exit__
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314__entry__
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Update/req
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Sample/req
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_final_index_sum_regn_update_start
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_scale_1/scale_rename_ack
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_complete/req
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_scale_1/scale_rename_req
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_scale_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/addr_of_1200_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_scale_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1238_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_resized_1
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1208_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1268_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_scaled_1
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1228_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_computed_1
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_resize_1/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/word_0/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_resize_1/$exit
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1218_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1258_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/ptr_deref_1204_Update/word_access_complete/word_0/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_resize_1/index_resize_ack
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/array_obj_ref_1199_index_resize_1/index_resize_req
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1278_Update/cr
      -- CP-element group 65: 	 branch_block_stmt_1090/assign_stmt_1201_to_assign_stmt_1314/type_cast_1248_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1090/merge_stmt_1186_PhiAck/$exit
      -- CP-element group 65: 	 branch_block_stmt_1090/merge_stmt_1186_PhiAck/phi_stmt_1187_ack
      -- 
    phi_stmt_1187_ack_3878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1187_ack_0, ack => sendOutput_CP_3266_elements(65)); -- 
    req_3515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => array_obj_ref_1199_index_offset_req_1); -- 
    req_3510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => array_obj_ref_1199_index_offset_req_0); -- 
    req_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => addr_of_1200_final_reg_req_1); -- 
    cr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1228_inst_req_1); -- 
    cr_3636_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3636_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1238_inst_req_1); -- 
    cr_3608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1218_inst_req_1); -- 
    cr_3664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1258_inst_req_1); -- 
    cr_3594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1208_inst_req_1); -- 
    cr_3678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1268_inst_req_1); -- 
    cr_3650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1248_inst_req_1); -- 
    cr_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => ptr_deref_1204_load_0_req_1); -- 
    cr_3692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => sendOutput_CP_3266_elements(65), ack => type_cast_1278_inst_req_1); -- 
    -- CP-element group 66:  merge  transition  place  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	58 
    -- CP-element group 66: 	9 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (16) 
      -- CP-element group 66: 	 branch_block_stmt_1090/branch_block_stmt_1090__exit__
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1325__exit__
      -- CP-element group 66: 	 branch_block_stmt_1090/return__
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1323__exit__
      -- CP-element group 66: 	 branch_block_stmt_1090/$exit
      -- CP-element group 66: 	 $exit
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1323_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1323_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1323_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1323_PhiAck/dummy
      -- CP-element group 66: 	 branch_block_stmt_1090/return___PhiReq/$entry
      -- CP-element group 66: 	 branch_block_stmt_1090/return___PhiReq/$exit
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1325_PhiReqMerge
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1325_PhiAck/$entry
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1325_PhiAck/$exit
      -- CP-element group 66: 	 branch_block_stmt_1090/merge_stmt_1325_PhiAck/dummy
      -- 
    sendOutput_CP_3266_elements(66) <= OrReduce(sendOutput_CP_3266_elements(58) & sendOutput_CP_3266_elements(9));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar_1198_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1198_scaled : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1199_root_address : std_logic_vector(13 downto 0);
    signal arrayidx_1201 : std_logic_vector(31 downto 0);
    signal cmp73_1142 : std_logic_vector(0 downto 0);
    signal conv17_1219 : std_logic_vector(7 downto 0);
    signal conv23_1229 : std_logic_vector(7 downto 0);
    signal conv29_1239 : std_logic_vector(7 downto 0);
    signal conv35_1249 : std_logic_vector(7 downto 0);
    signal conv41_1259 : std_logic_vector(7 downto 0);
    signal conv47_1269 : std_logic_vector(7 downto 0);
    signal conv53_1279 : std_logic_vector(7 downto 0);
    signal conv_1209 : std_logic_vector(7 downto 0);
    signal exitcond1_1314 : std_logic_vector(0 downto 0);
    signal iNsTr_0_1098 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1110 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1122 : std_logic_vector(31 downto 0);
    signal iNsTr_4_1171 : std_logic_vector(63 downto 0);
    signal indvar_1187 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1309 : std_logic_vector(63 downto 0);
    signal mul3_1136 : std_logic_vector(31 downto 0);
    signal mul_1131 : std_logic_vector(31 downto 0);
    signal ptr_deref_1101_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1101_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1101_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1101_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1101_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1113_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1113_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1113_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1113_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1113_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1125_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1125_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1125_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1125_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1125_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1204_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1204_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1204_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1204_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1204_word_offset_0 : std_logic_vector(13 downto 0);
    signal shr14_1215 : std_logic_vector(63 downto 0);
    signal shr20_1225 : std_logic_vector(63 downto 0);
    signal shr26_1235 : std_logic_vector(63 downto 0);
    signal shr32_1245 : std_logic_vector(63 downto 0);
    signal shr38_1255 : std_logic_vector(63 downto 0);
    signal shr44_1265 : std_logic_vector(63 downto 0);
    signal shr50_1275 : std_logic_vector(63 downto 0);
    signal tmp1_1114 : std_logic_vector(31 downto 0);
    signal tmp2_1126 : std_logic_vector(31 downto 0);
    signal tmp77_1155 : std_logic_vector(31 downto 0);
    signal tmp77x_xop_1167 : std_logic_vector(31 downto 0);
    signal tmp78_1161 : std_logic_vector(0 downto 0);
    signal tmp81_1184 : std_logic_vector(63 downto 0);
    signal tmp9_1205 : std_logic_vector(63 downto 0);
    signal tmp_1102 : std_logic_vector(31 downto 0);
    signal type_cast_1140_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1153_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1159_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1175_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1182_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1191_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1193_wire : std_logic_vector(63 downto 0);
    signal type_cast_1213_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1223_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1233_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1243_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1253_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1263_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1273_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1307_wire_constant : std_logic_vector(63 downto 0);
    signal xx_xop_1177 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    array_obj_ref_1199_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1199_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1199_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1199_resized_base_address <= "00000000000000";
    iNsTr_0_1098 <= "00000000000000000000000000000010";
    iNsTr_1_1110 <= "00000000000000000000000000000011";
    iNsTr_2_1122 <= "00000000000000000000000000000100";
    ptr_deref_1101_word_offset_0 <= "0000000";
    ptr_deref_1113_word_offset_0 <= "0000000";
    ptr_deref_1125_word_offset_0 <= "0000000";
    ptr_deref_1204_word_offset_0 <= "00000000000000";
    type_cast_1140_wire_constant <= "00000000000000000000000000000011";
    type_cast_1153_wire_constant <= "00000000000000000000000000000010";
    type_cast_1159_wire_constant <= "00000000000000000000000000000001";
    type_cast_1165_wire_constant <= "11111111111111111111111111111111";
    type_cast_1175_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1182_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1191_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1213_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1223_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1233_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1243_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1253_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1263_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1273_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1307_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    phi_stmt_1187: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1191_wire_constant & type_cast_1193_wire;
      req <= phi_stmt_1187_req_0 & phi_stmt_1187_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1187",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1187_ack_0,
          idata => idata,
          odata => indvar_1187,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1187
    -- flow-through select operator MUX_1183_inst
    tmp81_1184 <= xx_xop_1177 when (tmp78_1161(0) /=  '0') else type_cast_1182_wire_constant;
    addr_of_1200_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1200_final_reg_req_0;
      addr_of_1200_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1200_final_reg_req_1;
      addr_of_1200_final_reg_ack_1<= rack(0);
      addr_of_1200_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1200_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1199_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_1201,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1170_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1170_inst_req_0;
      type_cast_1170_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1170_inst_req_1;
      type_cast_1170_inst_ack_1<= rack(0);
      type_cast_1170_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1170_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp77x_xop_1167,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_4_1171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1193_inst_req_0;
      type_cast_1193_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1193_inst_req_1;
      type_cast_1193_inst_ack_1<= rack(0);
      type_cast_1193_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1193_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1309,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1193_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1208_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1208_inst_req_0;
      type_cast_1208_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1208_inst_req_1;
      type_cast_1208_inst_ack_1<= rack(0);
      type_cast_1208_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1208_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp9_1205,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_1209,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1218_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1218_inst_req_0;
      type_cast_1218_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1218_inst_req_1;
      type_cast_1218_inst_ack_1<= rack(0);
      type_cast_1218_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1218_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr14_1215,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv17_1219,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1228_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1228_inst_req_0;
      type_cast_1228_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1228_inst_req_1;
      type_cast_1228_inst_ack_1<= rack(0);
      type_cast_1228_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1228_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr20_1225,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv23_1229,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1238_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1238_inst_req_0;
      type_cast_1238_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1238_inst_req_1;
      type_cast_1238_inst_ack_1<= rack(0);
      type_cast_1238_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1238_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr26_1235,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv29_1239,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1248_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1248_inst_req_0;
      type_cast_1248_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1248_inst_req_1;
      type_cast_1248_inst_ack_1<= rack(0);
      type_cast_1248_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1248_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr32_1245,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv35_1249,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1258_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1258_inst_req_0;
      type_cast_1258_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1258_inst_req_1;
      type_cast_1258_inst_ack_1<= rack(0);
      type_cast_1258_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1258_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr38_1255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_1259,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1268_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1268_inst_req_0;
      type_cast_1268_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1268_inst_req_1;
      type_cast_1268_inst_ack_1<= rack(0);
      type_cast_1268_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1268_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr44_1265,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv47_1269,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1278_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1278_inst_req_0;
      type_cast_1278_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1278_inst_req_1;
      type_cast_1278_inst_ack_1<= rack(0);
      type_cast_1278_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1278_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => shr50_1275,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv53_1279,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1199_index_1_rename
    process(R_indvar_1198_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1198_resized;
      ov(13 downto 0) := iv;
      R_indvar_1198_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_index_1_resize
    process(indvar_1187) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1187;
      ov := iv(13 downto 0);
      R_indvar_1198_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1199_root_address_inst
    process(array_obj_ref_1199_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1199_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1199_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1101_addr_0
    process(ptr_deref_1101_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1101_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1101_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1101_base_resize
    process(iNsTr_0_1098) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_0_1098;
      ov := iv(6 downto 0);
      ptr_deref_1101_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1101_gather_scatter
    process(ptr_deref_1101_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1101_data_0;
      ov(31 downto 0) := iv;
      tmp_1102 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1101_root_address_inst
    process(ptr_deref_1101_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1101_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_addr_0
    process(ptr_deref_1113_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1113_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_base_resize
    process(iNsTr_1_1110) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_1110;
      ov := iv(6 downto 0);
      ptr_deref_1113_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_gather_scatter
    process(ptr_deref_1113_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_data_0;
      ov(31 downto 0) := iv;
      tmp1_1114 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1113_root_address_inst
    process(ptr_deref_1113_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1113_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1113_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_addr_0
    process(ptr_deref_1125_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_1125_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_base_resize
    process(iNsTr_2_1122) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_2_1122;
      ov := iv(6 downto 0);
      ptr_deref_1125_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_gather_scatter
    process(ptr_deref_1125_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_data_0;
      ov(31 downto 0) := iv;
      tmp2_1126 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1125_root_address_inst
    process(ptr_deref_1125_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1125_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_1125_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1204_addr_0
    process(ptr_deref_1204_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1204_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1204_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1204_base_resize
    process(arrayidx_1201) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_1201;
      ov := iv(13 downto 0);
      ptr_deref_1204_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1204_gather_scatter
    process(ptr_deref_1204_data_0) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1204_data_0;
      ov(63 downto 0) := iv;
      tmp9_1205 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1204_root_address_inst
    process(ptr_deref_1204_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1204_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1204_root_address <= ov(13 downto 0);
      --
    end process;
    if_stmt_1143_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp73_1142;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1143_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1143_branch_req_0,
          ack0 => if_stmt_1143_branch_ack_0,
          ack1 => if_stmt_1143_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1315_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_1314;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1315_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1315_branch_req_0,
          ack0 => if_stmt_1315_branch_ack_0,
          ack1 => if_stmt_1315_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1166_inst
    process(tmp77_1155) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp77_1155, type_cast_1165_wire_constant, tmp_var);
      tmp77x_xop_1167 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1176_inst
    process(iNsTr_4_1171) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_4_1171, type_cast_1175_wire_constant, tmp_var);
      xx_xop_1177 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1308_inst
    process(indvar_1187) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1187, type_cast_1307_wire_constant, tmp_var);
      indvarx_xnext_1309 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1313_inst
    process(indvarx_xnext_1309, tmp81_1184) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1309, tmp81_1184, tmp_var);
      exitcond1_1314 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1154_inst
    process(mul3_1136) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul3_1136, type_cast_1153_wire_constant, tmp_var);
      tmp77_1155 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1214_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1213_wire_constant, tmp_var);
      shr14_1215 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1224_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1223_wire_constant, tmp_var);
      shr20_1225 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1234_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1233_wire_constant, tmp_var);
      shr26_1235 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1244_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1243_wire_constant, tmp_var);
      shr32_1245 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1254_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1253_wire_constant, tmp_var);
      shr38_1255 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1264_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1263_wire_constant, tmp_var);
      shr44_1265 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_1274_inst
    process(tmp9_1205) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp9_1205, type_cast_1273_wire_constant, tmp_var);
      shr50_1275 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1130_inst
    process(tmp1_1114, tmp_1102) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp1_1114, tmp_1102, tmp_var);
      mul_1131 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_1135_inst
    process(mul_1131, tmp2_1126) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_1131, tmp2_1126, tmp_var);
      mul3_1136 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1141_inst
    process(mul3_1136) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul3_1136, type_cast_1140_wire_constant, tmp_var);
      cmp73_1142 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1160_inst
    process(tmp77_1155) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp77_1155, type_cast_1159_wire_constant, tmp_var);
      tmp78_1161 <= tmp_var; --
    end process;
    -- shared split operator group (16) : array_obj_ref_1199_index_offset 
    ApIntAdd_group_16: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1198_scaled;
      array_obj_ref_1199_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1199_index_offset_req_0;
      array_obj_ref_1199_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1199_index_offset_req_1;
      array_obj_ref_1199_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_16_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_16_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_16",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared load operator group (0) : ptr_deref_1101_load_0 ptr_deref_1113_load_0 ptr_deref_1125_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_1101_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1113_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1125_load_0_req_0;
      ptr_deref_1101_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1113_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1125_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1101_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1113_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1125_load_0_req_1;
      ptr_deref_1101_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1113_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1125_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1101_word_address_0 & ptr_deref_1113_word_address_0 & ptr_deref_1125_word_address_0;
      ptr_deref_1101_data_0 <= data_out(95 downto 64);
      ptr_deref_1113_data_0 <= data_out(63 downto 32);
      ptr_deref_1125_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1204_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1204_load_0_req_0;
      ptr_deref_1204_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1204_load_0_req_1;
      ptr_deref_1204_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1204_word_address_0;
      ptr_deref_1204_data_0 <= data_out(63 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 14,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(13 downto 0),
          mtag => memory_space_5_lr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(63 downto 0),
          mtag => memory_space_5_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared outport operator group (0) : WPIPE_ConvTranspose_output_pipe_1298_inst WPIPE_ConvTranspose_output_pipe_1286_inst WPIPE_ConvTranspose_output_pipe_1295_inst WPIPE_ConvTranspose_output_pipe_1292_inst WPIPE_ConvTranspose_output_pipe_1283_inst WPIPE_ConvTranspose_output_pipe_1289_inst WPIPE_ConvTranspose_output_pipe_1280_inst WPIPE_ConvTranspose_output_pipe_1301_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal sample_req, sample_ack : BooleanArray( 7 downto 0);
      signal update_req, update_ack : BooleanArray( 7 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 7 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      constant inBUFs : IntegerArray(7 downto 0) := (7 => 0, 6 => 0, 5 => 0, 4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(7 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false);
      constant guardBuffering: IntegerArray(7 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2);
      -- 
    begin -- 
      sample_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_0;
      sample_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_0;
      sample_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_0;
      sample_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_0;
      sample_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_0;
      sample_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_0;
      sample_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_0;
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_0 <= sample_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_0 <= sample_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_0 <= sample_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_0 <= sample_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_0 <= sample_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_0 <= sample_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(7) <= WPIPE_ConvTranspose_output_pipe_1298_inst_req_1;
      update_req_unguarded(6) <= WPIPE_ConvTranspose_output_pipe_1286_inst_req_1;
      update_req_unguarded(5) <= WPIPE_ConvTranspose_output_pipe_1295_inst_req_1;
      update_req_unguarded(4) <= WPIPE_ConvTranspose_output_pipe_1292_inst_req_1;
      update_req_unguarded(3) <= WPIPE_ConvTranspose_output_pipe_1283_inst_req_1;
      update_req_unguarded(2) <= WPIPE_ConvTranspose_output_pipe_1289_inst_req_1;
      update_req_unguarded(1) <= WPIPE_ConvTranspose_output_pipe_1280_inst_req_1;
      update_req_unguarded(0) <= WPIPE_ConvTranspose_output_pipe_1301_inst_req_1;
      WPIPE_ConvTranspose_output_pipe_1298_inst_ack_1 <= update_ack_unguarded(7);
      WPIPE_ConvTranspose_output_pipe_1286_inst_ack_1 <= update_ack_unguarded(6);
      WPIPE_ConvTranspose_output_pipe_1295_inst_ack_1 <= update_ack_unguarded(5);
      WPIPE_ConvTranspose_output_pipe_1292_inst_ack_1 <= update_ack_unguarded(4);
      WPIPE_ConvTranspose_output_pipe_1283_inst_ack_1 <= update_ack_unguarded(3);
      WPIPE_ConvTranspose_output_pipe_1289_inst_ack_1 <= update_ack_unguarded(2);
      WPIPE_ConvTranspose_output_pipe_1280_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_ConvTranspose_output_pipe_1301_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      data_in <= conv17_1219 & conv41_1259 & conv23_1229 & conv29_1239 & conv47_1269 & conv35_1249 & conv53_1279 & conv_1209;
      ConvTranspose_output_pipe_write_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_output_pipe_write_0_gI", nreqs => 8, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_output_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "ConvTranspose_output_pipe", data_width => 8, num_reqs => 8, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => ConvTranspose_output_pipe_pipe_write_req(0),
          oack => ConvTranspose_output_pipe_pipe_write_ack(0),
          odata => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end sendOutput_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity testConfigure is -- 
  generic (tag_length : integer); 
  port ( -- 
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
    memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
    memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity testConfigure;
architecture testConfigure_arch of testConfigure is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 16)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ret_val_x_x_update_enable: Boolean;
  signal testConfigure_CP_0_start: Boolean;
  signal testConfigure_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal RPIPE_ConvTranspose_input_pipe_874_inst_req_1 : boolean;
  signal type_cast_896_inst_req_1 : boolean;
  signal ptr_deref_467_load_0_ack_1 : boolean;
  signal if_stmt_936_branch_ack_0 : boolean;
  signal ptr_deref_381_load_0_req_0 : boolean;
  signal addr_of_1054_final_reg_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_req_0 : boolean;
  signal if_stmt_500_branch_ack_1 : boolean;
  signal if_stmt_500_branch_ack_0 : boolean;
  signal array_obj_ref_1053_index_offset_ack_0 : boolean;
  signal if_stmt_500_branch_req_0 : boolean;
  signal ptr_deref_381_load_0_ack_0 : boolean;
  signal type_cast_38_inst_req_0 : boolean;
  signal type_cast_38_inst_ack_0 : boolean;
  signal ptr_deref_368_store_0_ack_1 : boolean;
  signal ptr_deref_368_store_0_req_1 : boolean;
  signal type_cast_357_inst_req_0 : boolean;
  signal ptr_deref_368_store_0_ack_0 : boolean;
  signal ptr_deref_368_store_0_req_0 : boolean;
  signal type_cast_357_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 : boolean;
  signal ptr_deref_467_load_0_req_1 : boolean;
  signal type_cast_38_inst_req_1 : boolean;
  signal type_cast_38_inst_ack_1 : boolean;
  signal ptr_deref_47_store_0_req_0 : boolean;
  signal ptr_deref_47_store_0_ack_0 : boolean;
  signal ptr_deref_47_store_0_req_1 : boolean;
  signal ptr_deref_47_store_0_ack_1 : boolean;
  signal type_cast_357_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_874_inst_ack_1 : boolean;
  signal type_cast_62_inst_req_0 : boolean;
  signal type_cast_62_inst_ack_0 : boolean;
  signal type_cast_62_inst_req_1 : boolean;
  signal type_cast_62_inst_ack_1 : boolean;
  signal if_stmt_64_branch_req_0 : boolean;
  signal if_stmt_64_branch_ack_1 : boolean;
  signal if_stmt_64_branch_ack_0 : boolean;
  signal type_cast_95_inst_req_0 : boolean;
  signal type_cast_95_inst_ack_0 : boolean;
  signal array_obj_ref_1053_index_offset_req_1 : boolean;
  signal type_cast_95_inst_req_1 : boolean;
  signal type_cast_95_inst_ack_1 : boolean;
  signal array_obj_ref_101_index_offset_req_0 : boolean;
  signal array_obj_ref_101_index_offset_ack_0 : boolean;
  signal array_obj_ref_101_index_offset_req_1 : boolean;
  signal array_obj_ref_101_index_offset_ack_1 : boolean;
  signal ptr_deref_467_load_0_ack_0 : boolean;
  signal ptr_deref_455_load_0_ack_1 : boolean;
  signal addr_of_102_final_reg_req_0 : boolean;
  signal addr_of_102_final_reg_ack_0 : boolean;
  signal addr_of_102_final_reg_req_1 : boolean;
  signal ptr_deref_979_load_0_req_1 : boolean;
  signal addr_of_102_final_reg_ack_1 : boolean;
  signal type_cast_486_inst_ack_1 : boolean;
  signal type_cast_914_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_req_1 : boolean;
  signal ptr_deref_431_load_0_ack_1 : boolean;
  signal ptr_deref_431_load_0_req_1 : boolean;
  signal ptr_deref_455_load_0_req_1 : boolean;
  signal type_cast_896_inst_ack_1 : boolean;
  signal ptr_deref_105_store_0_req_0 : boolean;
  signal ptr_deref_105_store_0_ack_0 : boolean;
  signal ptr_deref_105_store_0_req_1 : boolean;
  signal ptr_deref_105_store_0_ack_1 : boolean;
  signal if_stmt_997_branch_ack_0 : boolean;
  signal type_cast_486_inst_req_1 : boolean;
  signal ptr_deref_979_load_0_ack_0 : boolean;
  signal addr_of_274_final_reg_req_0 : boolean;
  signal type_cast_878_inst_req_1 : boolean;
  signal addr_of_274_final_reg_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_ack_0 : boolean;
  signal addr_of_274_final_reg_req_1 : boolean;
  signal addr_of_274_final_reg_ack_1 : boolean;
  signal ptr_deref_393_load_0_ack_1 : boolean;
  signal ptr_deref_393_load_0_req_1 : boolean;
  signal type_cast_914_inst_req_0 : boolean;
  signal ptr_deref_405_load_0_ack_1 : boolean;
  signal ptr_deref_122_load_0_req_0 : boolean;
  signal ptr_deref_122_load_0_ack_0 : boolean;
  signal ptr_deref_122_load_0_req_1 : boolean;
  signal ptr_deref_122_load_0_ack_1 : boolean;
  signal ptr_deref_443_load_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_130_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_req_0 : boolean;
  signal type_cast_134_inst_req_0 : boolean;
  signal type_cast_134_inst_ack_0 : boolean;
  signal ptr_deref_443_load_0_req_1 : boolean;
  signal type_cast_134_inst_req_1 : boolean;
  signal type_cast_134_inst_ack_1 : boolean;
  signal addr_of_1054_final_reg_ack_1 : boolean;
  signal ptr_deref_467_load_0_req_0 : boolean;
  signal ptr_deref_405_load_0_req_1 : boolean;
  signal if_stmt_136_branch_req_0 : boolean;
  signal if_stmt_136_branch_ack_1 : boolean;
  signal if_stmt_136_branch_ack_0 : boolean;
  signal ptr_deref_431_load_0_ack_0 : boolean;
  signal ptr_deref_431_load_0_req_0 : boolean;
  signal type_cast_419_inst_ack_1 : boolean;
  signal ptr_deref_164_store_0_req_0 : boolean;
  signal ptr_deref_164_store_0_ack_0 : boolean;
  signal ptr_deref_455_load_0_ack_0 : boolean;
  signal ptr_deref_164_store_0_req_1 : boolean;
  signal ptr_deref_164_store_0_ack_1 : boolean;
  signal type_cast_486_inst_ack_0 : boolean;
  signal type_cast_357_inst_ack_0 : boolean;
  signal if_stmt_173_branch_req_0 : boolean;
  signal if_stmt_173_branch_ack_1 : boolean;
  signal if_stmt_173_branch_ack_0 : boolean;
  signal type_cast_419_inst_req_1 : boolean;
  signal type_cast_198_inst_req_0 : boolean;
  signal ptr_deref_979_load_0_ack_1 : boolean;
  signal type_cast_198_inst_ack_0 : boolean;
  signal ptr_deref_443_load_0_ack_0 : boolean;
  signal type_cast_198_inst_req_1 : boolean;
  signal type_cast_198_inst_ack_1 : boolean;
  signal type_cast_486_inst_req_0 : boolean;
  signal ptr_deref_455_load_0_req_0 : boolean;
  signal array_obj_ref_204_index_offset_req_0 : boolean;
  signal array_obj_ref_204_index_offset_ack_0 : boolean;
  signal array_obj_ref_204_index_offset_req_1 : boolean;
  signal array_obj_ref_204_index_offset_ack_1 : boolean;
  signal type_cast_419_inst_ack_0 : boolean;
  signal addr_of_205_final_reg_req_0 : boolean;
  signal addr_of_205_final_reg_ack_0 : boolean;
  signal ptr_deref_405_load_0_ack_0 : boolean;
  signal ptr_deref_443_load_0_req_0 : boolean;
  signal addr_of_205_final_reg_req_1 : boolean;
  signal type_cast_419_inst_req_0 : boolean;
  signal addr_of_205_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_208_inst_ack_1 : boolean;
  signal type_cast_212_inst_req_0 : boolean;
  signal type_cast_212_inst_ack_0 : boolean;
  signal type_cast_212_inst_req_1 : boolean;
  signal type_cast_212_inst_ack_1 : boolean;
  signal ptr_deref_215_store_0_req_0 : boolean;
  signal ptr_deref_215_store_0_ack_0 : boolean;
  signal ptr_deref_215_store_0_req_1 : boolean;
  signal ptr_deref_215_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_856_inst_ack_1 : boolean;
  signal ptr_deref_405_load_0_req_0 : boolean;
  signal ptr_deref_381_load_0_ack_1 : boolean;
  signal ptr_deref_232_load_0_req_0 : boolean;
  signal ptr_deref_232_load_0_ack_0 : boolean;
  signal ptr_deref_381_load_0_req_1 : boolean;
  signal ptr_deref_232_load_0_req_1 : boolean;
  signal ptr_deref_232_load_0_ack_1 : boolean;
  signal if_stmt_239_branch_req_0 : boolean;
  signal if_stmt_239_branch_ack_1 : boolean;
  signal if_stmt_239_branch_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_249_inst_ack_1 : boolean;
  signal type_cast_253_inst_req_0 : boolean;
  signal type_cast_253_inst_ack_0 : boolean;
  signal type_cast_253_inst_req_1 : boolean;
  signal type_cast_253_inst_ack_1 : boolean;
  signal array_obj_ref_1053_index_offset_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_ack_0 : boolean;
  signal ptr_deref_277_store_0_req_0 : boolean;
  signal ptr_deref_277_store_0_ack_0 : boolean;
  signal ptr_deref_277_store_0_req_1 : boolean;
  signal ptr_deref_277_store_0_ack_1 : boolean;
  signal type_cast_914_inst_req_1 : boolean;
  signal ptr_deref_393_load_0_ack_0 : boolean;
  signal ptr_deref_393_load_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 : boolean;
  signal ptr_deref_955_load_0_req_0 : boolean;
  signal type_cast_285_inst_req_0 : boolean;
  signal type_cast_285_inst_ack_0 : boolean;
  signal type_cast_285_inst_req_1 : boolean;
  signal type_cast_285_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_req_1 : boolean;
  signal type_cast_878_inst_req_0 : boolean;
  signal if_stmt_299_branch_req_0 : boolean;
  signal type_cast_914_inst_ack_1 : boolean;
  signal if_stmt_299_branch_ack_1 : boolean;
  signal if_stmt_299_branch_ack_0 : boolean;
  signal type_cast_878_inst_ack_0 : boolean;
  signal STORE_padding_311_store_0_req_0 : boolean;
  signal STORE_padding_311_store_0_ack_0 : boolean;
  signal STORE_padding_311_store_0_req_1 : boolean;
  signal ptr_deref_955_load_0_ack_0 : boolean;
  signal STORE_padding_311_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_315_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_910_inst_ack_1 : boolean;
  signal type_cast_319_inst_req_0 : boolean;
  signal type_cast_319_inst_ack_0 : boolean;
  signal type_cast_319_inst_req_1 : boolean;
  signal type_cast_319_inst_ack_1 : boolean;
  signal type_cast_860_inst_req_0 : boolean;
  signal type_cast_860_inst_ack_0 : boolean;
  signal ptr_deref_330_store_0_req_0 : boolean;
  signal ptr_deref_330_store_0_ack_0 : boolean;
  signal ptr_deref_330_store_0_req_1 : boolean;
  signal ptr_deref_330_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_334_inst_ack_1 : boolean;
  signal type_cast_338_inst_req_0 : boolean;
  signal type_cast_338_inst_ack_0 : boolean;
  signal type_cast_338_inst_req_1 : boolean;
  signal type_cast_338_inst_ack_1 : boolean;
  signal ptr_deref_349_store_0_req_0 : boolean;
  signal ptr_deref_349_store_0_ack_0 : boolean;
  signal ptr_deref_349_store_0_req_1 : boolean;
  signal ptr_deref_349_store_0_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 : boolean;
  signal array_obj_ref_1053_index_offset_req_0 : boolean;
  signal if_stmt_521_branch_req_0 : boolean;
  signal if_stmt_936_branch_ack_1 : boolean;
  signal if_stmt_521_branch_ack_1 : boolean;
  signal if_stmt_521_branch_ack_0 : boolean;
  signal type_cast_860_inst_ack_1 : boolean;
  signal type_cast_860_inst_req_1 : boolean;
  signal ptr_deref_979_load_0_req_0 : boolean;
  signal if_stmt_997_branch_ack_1 : boolean;
  signal type_cast_540_inst_req_0 : boolean;
  signal type_cast_540_inst_ack_0 : boolean;
  signal type_cast_540_inst_req_1 : boolean;
  signal type_cast_540_inst_ack_1 : boolean;
  signal addr_of_1054_final_reg_ack_0 : boolean;
  signal if_stmt_936_branch_req_0 : boolean;
  signal array_obj_ref_575_index_offset_req_0 : boolean;
  signal array_obj_ref_575_index_offset_ack_0 : boolean;
  signal array_obj_ref_575_index_offset_req_1 : boolean;
  signal array_obj_ref_575_index_offset_ack_1 : boolean;
  signal addr_of_1054_final_reg_req_0 : boolean;
  signal type_cast_896_inst_ack_0 : boolean;
  signal addr_of_576_final_reg_req_0 : boolean;
  signal addr_of_576_final_reg_ack_0 : boolean;
  signal addr_of_576_final_reg_req_1 : boolean;
  signal addr_of_576_final_reg_ack_1 : boolean;
  signal type_cast_896_inst_req_0 : boolean;
  signal ptr_deref_922_store_0_ack_1 : boolean;
  signal ptr_deref_922_store_0_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 : boolean;
  signal type_cast_583_inst_req_0 : boolean;
  signal type_cast_583_inst_ack_0 : boolean;
  signal type_cast_583_inst_req_1 : boolean;
  signal type_cast_583_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_592_inst_ack_1 : boolean;
  signal if_stmt_997_branch_req_0 : boolean;
  signal type_cast_596_inst_req_0 : boolean;
  signal type_cast_596_inst_ack_0 : boolean;
  signal type_cast_596_inst_req_1 : boolean;
  signal type_cast_596_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_610_inst_ack_1 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal type_cast_614_inst_req_1 : boolean;
  signal type_cast_614_inst_ack_1 : boolean;
  signal ptr_deref_1057_store_0_ack_0 : boolean;
  signal type_cast_1024_inst_ack_1 : boolean;
  signal type_cast_1024_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_628_inst_ack_1 : boolean;
  signal type_cast_632_inst_req_0 : boolean;
  signal type_cast_632_inst_ack_0 : boolean;
  signal type_cast_632_inst_req_1 : boolean;
  signal type_cast_632_inst_ack_1 : boolean;
  signal ptr_deref_1057_store_0_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_646_inst_ack_1 : boolean;
  signal ptr_deref_922_store_0_ack_0 : boolean;
  signal ptr_deref_922_store_0_req_0 : boolean;
  signal type_cast_650_inst_req_0 : boolean;
  signal type_cast_650_inst_ack_0 : boolean;
  signal type_cast_650_inst_req_1 : boolean;
  signal type_cast_650_inst_ack_1 : boolean;
  signal type_cast_1024_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 : boolean;
  signal type_cast_668_inst_req_0 : boolean;
  signal ptr_deref_967_load_0_ack_1 : boolean;
  signal type_cast_668_inst_ack_0 : boolean;
  signal type_cast_668_inst_req_1 : boolean;
  signal ptr_deref_967_load_0_req_1 : boolean;
  signal type_cast_668_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_892_inst_req_0 : boolean;
  signal type_cast_1024_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 : boolean;
  signal type_cast_686_inst_req_0 : boolean;
  signal type_cast_686_inst_ack_0 : boolean;
  signal type_cast_686_inst_req_1 : boolean;
  signal type_cast_686_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 : boolean;
  signal type_cast_704_inst_req_0 : boolean;
  signal ptr_deref_967_load_0_ack_0 : boolean;
  signal type_cast_704_inst_ack_0 : boolean;
  signal type_cast_704_inst_req_1 : boolean;
  signal ptr_deref_967_load_0_req_0 : boolean;
  signal type_cast_704_inst_ack_1 : boolean;
  signal ptr_deref_712_store_0_req_0 : boolean;
  signal ptr_deref_712_store_0_ack_0 : boolean;
  signal type_cast_842_inst_ack_1 : boolean;
  signal ptr_deref_712_store_0_req_1 : boolean;
  signal ptr_deref_712_store_0_ack_1 : boolean;
  signal type_cast_842_inst_req_1 : boolean;
  signal ptr_deref_955_load_0_ack_1 : boolean;
  signal if_stmt_726_branch_req_0 : boolean;
  signal ptr_deref_955_load_0_req_1 : boolean;
  signal if_stmt_726_branch_ack_1 : boolean;
  signal if_stmt_726_branch_ack_0 : boolean;
  signal type_cast_750_inst_req_0 : boolean;
  signal type_cast_750_inst_ack_0 : boolean;
  signal type_cast_750_inst_req_1 : boolean;
  signal type_cast_750_inst_ack_1 : boolean;
  signal type_cast_878_inst_ack_1 : boolean;
  signal array_obj_ref_785_index_offset_req_0 : boolean;
  signal array_obj_ref_785_index_offset_ack_0 : boolean;
  signal array_obj_ref_785_index_offset_req_1 : boolean;
  signal array_obj_ref_785_index_offset_ack_1 : boolean;
  signal addr_of_786_final_reg_req_0 : boolean;
  signal addr_of_786_final_reg_ack_0 : boolean;
  signal addr_of_786_final_reg_req_1 : boolean;
  signal addr_of_786_final_reg_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 : boolean;
  signal type_cast_793_inst_req_0 : boolean;
  signal type_cast_793_inst_ack_0 : boolean;
  signal type_cast_793_inst_req_1 : boolean;
  signal type_cast_793_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_802_inst_ack_1 : boolean;
  signal type_cast_806_inst_req_0 : boolean;
  signal type_cast_806_inst_ack_0 : boolean;
  signal type_cast_806_inst_req_1 : boolean;
  signal type_cast_806_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_820_inst_ack_1 : boolean;
  signal type_cast_824_inst_req_0 : boolean;
  signal type_cast_824_inst_ack_0 : boolean;
  signal type_cast_824_inst_req_1 : boolean;
  signal type_cast_824_inst_ack_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_req_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_ack_0 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_req_1 : boolean;
  signal RPIPE_ConvTranspose_input_pipe_838_inst_ack_1 : boolean;
  signal type_cast_842_inst_req_0 : boolean;
  signal type_cast_842_inst_ack_0 : boolean;
  signal ptr_deref_1057_store_0_req_1 : boolean;
  signal ptr_deref_1057_store_0_ack_1 : boolean;
  signal if_stmt_1072_branch_req_0 : boolean;
  signal if_stmt_1072_branch_ack_1 : boolean;
  signal if_stmt_1072_branch_ack_0 : boolean;
  signal type_cast_1083_inst_req_0 : boolean;
  signal type_cast_1083_inst_ack_0 : boolean;
  signal type_cast_1083_inst_req_1 : boolean;
  signal type_cast_1083_inst_ack_1 : boolean;
  signal type_cast_76_inst_req_0 : boolean;
  signal type_cast_76_inst_ack_0 : boolean;
  signal type_cast_76_inst_req_1 : boolean;
  signal type_cast_76_inst_ack_1 : boolean;
  signal phi_stmt_73_req_0 : boolean;
  signal type_cast_83_inst_req_0 : boolean;
  signal type_cast_83_inst_ack_0 : boolean;
  signal type_cast_83_inst_req_1 : boolean;
  signal type_cast_83_inst_ack_1 : boolean;
  signal phi_stmt_80_req_0 : boolean;
  signal phi_stmt_73_req_1 : boolean;
  signal type_cast_85_inst_req_0 : boolean;
  signal type_cast_85_inst_ack_0 : boolean;
  signal type_cast_85_inst_req_1 : boolean;
  signal type_cast_85_inst_ack_1 : boolean;
  signal phi_stmt_80_req_1 : boolean;
  signal phi_stmt_73_ack_0 : boolean;
  signal phi_stmt_80_ack_0 : boolean;
  signal type_cast_146_inst_req_0 : boolean;
  signal type_cast_146_inst_ack_0 : boolean;
  signal type_cast_146_inst_req_1 : boolean;
  signal type_cast_146_inst_ack_1 : boolean;
  signal phi_stmt_143_req_0 : boolean;
  signal phi_stmt_143_ack_0 : boolean;
  signal type_cast_153_inst_req_0 : boolean;
  signal type_cast_153_inst_ack_0 : boolean;
  signal type_cast_153_inst_req_1 : boolean;
  signal type_cast_153_inst_ack_1 : boolean;
  signal phi_stmt_150_req_0 : boolean;
  signal type_cast_155_inst_req_0 : boolean;
  signal type_cast_155_inst_ack_0 : boolean;
  signal type_cast_155_inst_req_1 : boolean;
  signal type_cast_155_inst_ack_1 : boolean;
  signal phi_stmt_150_req_1 : boolean;
  signal phi_stmt_150_ack_0 : boolean;
  signal type_cast_185_inst_req_0 : boolean;
  signal type_cast_185_inst_ack_0 : boolean;
  signal type_cast_185_inst_req_1 : boolean;
  signal type_cast_185_inst_ack_1 : boolean;
  signal phi_stmt_182_req_0 : boolean;
  signal phi_stmt_182_req_1 : boolean;
  signal phi_stmt_182_ack_0 : boolean;
  signal phi_stmt_257_req_0 : boolean;
  signal type_cast_267_inst_req_0 : boolean;
  signal type_cast_267_inst_ack_0 : boolean;
  signal type_cast_267_inst_req_1 : boolean;
  signal type_cast_267_inst_ack_1 : boolean;
  signal phi_stmt_264_req_0 : boolean;
  signal type_cast_263_inst_req_0 : boolean;
  signal type_cast_263_inst_ack_0 : boolean;
  signal type_cast_263_inst_req_1 : boolean;
  signal type_cast_263_inst_ack_1 : boolean;
  signal phi_stmt_257_req_1 : boolean;
  signal type_cast_269_inst_req_0 : boolean;
  signal type_cast_269_inst_ack_0 : boolean;
  signal type_cast_269_inst_req_1 : boolean;
  signal type_cast_269_inst_ack_1 : boolean;
  signal phi_stmt_264_req_1 : boolean;
  signal phi_stmt_257_ack_0 : boolean;
  signal phi_stmt_264_ack_0 : boolean;
  signal type_cast_309_inst_req_0 : boolean;
  signal type_cast_309_inst_ack_0 : boolean;
  signal type_cast_309_inst_req_1 : boolean;
  signal type_cast_309_inst_ack_1 : boolean;
  signal phi_stmt_306_req_0 : boolean;
  signal phi_stmt_306_ack_0 : boolean;
  signal phi_stmt_563_req_0 : boolean;
  signal type_cast_569_inst_req_0 : boolean;
  signal type_cast_569_inst_ack_0 : boolean;
  signal type_cast_569_inst_req_1 : boolean;
  signal type_cast_569_inst_ack_1 : boolean;
  signal phi_stmt_563_req_1 : boolean;
  signal phi_stmt_563_ack_0 : boolean;
  signal phi_stmt_773_req_0 : boolean;
  signal type_cast_779_inst_req_0 : boolean;
  signal type_cast_779_inst_ack_0 : boolean;
  signal type_cast_779_inst_req_1 : boolean;
  signal type_cast_779_inst_ack_1 : boolean;
  signal phi_stmt_773_req_1 : boolean;
  signal phi_stmt_773_ack_0 : boolean;
  signal phi_stmt_1041_req_0 : boolean;
  signal type_cast_1047_inst_req_0 : boolean;
  signal type_cast_1047_inst_ack_0 : boolean;
  signal type_cast_1047_inst_req_1 : boolean;
  signal type_cast_1047_inst_ack_1 : boolean;
  signal phi_stmt_1041_req_1 : boolean;
  signal phi_stmt_1041_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "testConfigure_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  testConfigure_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "testConfigure_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 16) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(15 downto 0) <= ret_val_x_x_buffer;
  ret_val_x_x <= out_buffer_data_out(15 downto 0);
  out_buffer_data_in(tag_length + 15 downto 16) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 15 downto 16);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= testConfigure_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  testConfigure_CP_0: Block -- control-path 
    signal testConfigure_CP_0_elements: BooleanArray(310 downto 0);
    -- 
  begin -- 
    testConfigure_CP_0_elements(0) <= testConfigure_CP_0_start;
    testConfigure_CP_0_symbol <= testConfigure_CP_0_elements(233);
    -- CP-element group 0:  fork  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	5 
    -- CP-element group 0: 	7 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (35) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_32/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/branch_block_stmt_32__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__entry__
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/rr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_root_address_calculated
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_address_resized
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_addr_resize/base_resize_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/$exit
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_req
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_word_addrgen/root_register_ack
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/cr
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_start_
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$entry
      -- CP-element group 0: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/cr
      -- 
    rr_118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_0); -- 
    cr_137_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_137_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_38_inst_req_1); -- 
    cr_187_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_187_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => ptr_deref_47_store_0_req_1); -- 
    cr_215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(0), ack => type_cast_62_inst_req_1); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_start_
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Sample/ra
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/cr
      -- 
    ra_119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_0, ack => testConfigure_CP_0_elements(1)); -- 
    cr_123_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_123_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(1), ack => RPIPE_ConvTranspose_input_pipe_34_inst_req_1); -- 
    -- CP-element group 2:  fork  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (9) 
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/rr
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_34_Update/ca
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/rr
      -- 
    ca_124_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_34_inst_ack_1, ack => testConfigure_CP_0_elements(2)); -- 
    rr_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => type_cast_38_inst_req_0); -- 
    rr_196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(2), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Sample/ra
      -- CP-element group 3: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_sample_completed_
      -- 
    ra_133_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_0, ack => testConfigure_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_38_Update/ca
      -- 
    ca_138_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_38_inst_ack_1, ack => testConfigure_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (9) 
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/$exit
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_req
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/ptr_deref_47_Split/split_ack
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$entry
      -- CP-element group 5: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/rr
      -- 
    rr_176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(5), ack => ptr_deref_47_store_0_req_0); -- 
    testConfigure_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "testConfigure_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(0) & testConfigure_CP_0_elements(4);
      gj_testConfigure_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_sample_completed_
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/$exit
      -- CP-element group 6: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Sample/word_access_start/word_0/ra
      -- 
    ra_177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_0, ack => testConfigure_CP_0_elements(6)); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	0 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (5) 
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_update_completed_
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/$exit
      -- CP-element group 7: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/ptr_deref_47_Update/word_access_complete/word_0/ca
      -- 
    ca_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_47_store_0_ack_1, ack => testConfigure_CP_0_elements(7)); -- 
    -- CP-element group 8:  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_start_
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Sample/ra
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/cr
      -- 
    ra_197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_0, ack => testConfigure_CP_0_elements(8)); -- 
    cr_201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(8), ack => RPIPE_ConvTranspose_input_pipe_58_inst_req_1); -- 
    -- CP-element group 9:  transition  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9:  members (6) 
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/RPIPE_ConvTranspose_input_pipe_58_Update/ca
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_start_
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/rr
      -- 
    ca_202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_58_inst_ack_1, ack => testConfigure_CP_0_elements(9)); -- 
    rr_210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(9), ack => type_cast_62_inst_req_0); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Sample/ra
      -- 
    ra_211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_0, ack => testConfigure_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/type_cast_62_Update/ca
      -- 
    ca_216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_62_inst_ack_1, ack => testConfigure_CP_0_elements(11)); -- 
    -- CP-element group 12:  branch  join  transition  place  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (10) 
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63__exit__
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64__entry__
      -- CP-element group 12: 	 branch_block_stmt_32/assign_stmt_35_to_assign_stmt_63/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_dead_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/$exit
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_eval_test/branch_req
      -- CP-element group 12: 	 branch_block_stmt_32/R_cmp227_65_place
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_if_link/$entry
      -- CP-element group 12: 	 branch_block_stmt_32/if_stmt_64_else_link/$entry
      -- 
    branch_req_224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(12), ack => if_stmt_64_branch_req_0); -- 
    testConfigure_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(7) & testConfigure_CP_0_elements(11);
      gj_testConfigure_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  fork  transition  place  input  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	254 
    -- CP-element group 13: 	255 
    -- CP-element group 13:  members (12) 
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/$exit
      -- CP-element group 13: 	 branch_block_stmt_32/if_stmt_64_if_link/if_choice_transition
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/rr
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$entry
      -- CP-element group 13: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/cr
      -- 
    if_choice_transition_229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_1, ack => testConfigure_CP_0_elements(13)); -- 
    rr_2787_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2787_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_153_inst_req_0); -- 
    cr_2792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(13), ack => type_cast_153_inst_req_1); -- 
    -- CP-element group 14:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	241 
    -- CP-element group 14: 	242 
    -- CP-element group 14: 	243 
    -- CP-element group 14:  members (22) 
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70__exit__
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/if_stmt_64_else_link/else_choice_transition
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/entry_forx_xbodyx_xpreheader_PhiReq/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiReqMerge
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/$exit
      -- CP-element group 14: 	 branch_block_stmt_32/merge_stmt_70_PhiAck/dummy
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/cr
      -- 
    else_choice_transition_233_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_64_branch_ack_0, ack => testConfigure_CP_0_elements(14)); -- 
    rr_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_0); -- 
    cr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(14), ack => type_cast_85_inst_req_1); -- 
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	249 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/ra
      -- 
    ra_247_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_0, ack => testConfigure_CP_0_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	249 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	31 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/ca
      -- 
    ca_252_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_95_inst_ack_1, ack => testConfigure_CP_0_elements(16)); -- 
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	249 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	31 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_sample_complete
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/$exit
      -- CP-element group 17: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/ack
      -- 
    ack_278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_0, ack => testConfigure_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	249 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (11) 
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_root_address_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_offset_calculated
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/$exit
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/sum_rename_req
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_base_plus_offset/sum_rename_ack
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/$entry
      -- CP-element group 18: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/req
      -- 
    ack_283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_101_index_offset_ack_1, ack => testConfigure_CP_0_elements(18)); -- 
    req_292_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_292_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(18), ack => addr_of_102_final_reg_req_0); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/$exit
      -- CP-element group 19: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_request/ack
      -- 
    ack_293_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_0, ack => testConfigure_CP_0_elements(19)); -- 
    -- CP-element group 20:  join  fork  transition  input  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	249 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (28) 
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_sample_start_
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_root_address_calculated
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_address_resized
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/base_resize_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_addr_resize/base_resize_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/sum_rename_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_base_plus_offset/sum_rename_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/root_register_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_word_addrgen/root_register_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/$exit
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/split_req
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/ptr_deref_105_Split/split_ack
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/$entry
      -- CP-element group 20: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/rr
      -- 
    ack_298_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_102_final_reg_ack_1, ack => testConfigure_CP_0_elements(20)); -- 
    rr_336_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_336_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(20), ack => ptr_deref_105_store_0_req_0); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	30 
    -- CP-element group 21:  members (5) 
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_sample_completed_
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/$exit
      -- CP-element group 21: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Sample/word_access_start/word_0/ra
      -- 
    ra_337_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_0, ack => testConfigure_CP_0_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	249 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	31 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_update_completed_
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/$exit
      -- CP-element group 22: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/ca
      -- 
    ca_348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_105_store_0_ack_1, ack => testConfigure_CP_0_elements(22)); -- 
    -- CP-element group 23:  join  transition  output  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	30 
    -- CP-element group 23: 	249 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (5) 
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_sample_start_
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/$entry
      -- CP-element group 23: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/rr
      -- 
    rr_381_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_381_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(23), ack => ptr_deref_122_load_0_req_0); -- 
    testConfigure_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(30) & testConfigure_CP_0_elements(249);
      gj_testConfigure_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  transition  input  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (5) 
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_sample_completed_
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/$exit
      -- CP-element group 24: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Sample/word_access_start/word_0/ra
      -- 
    ra_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_0, ack => testConfigure_CP_0_elements(24)); -- 
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	249 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	31 
    -- CP-element group 25:  members (9) 
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/ca
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/$entry
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/$exit
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/merge_req
      -- CP-element group 25: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/ptr_deref_122_Merge/merge_ack
      -- 
    ca_393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_122_load_0_ack_1, ack => testConfigure_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	249 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_update_start_
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/ra
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/cr
      -- 
    ra_407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_130_inst_ack_0, ack => testConfigure_CP_0_elements(26)); -- 
    cr_411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(26), ack => RPIPE_ConvTranspose_input_pipe_130_inst_req_1); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Update/ca
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/$entry
      -- CP-element group 27: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/rr
      -- 
    ca_412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_130_inst_ack_1, ack => testConfigure_CP_0_elements(27)); -- 
    rr_420_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_420_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(27), ack => type_cast_134_inst_req_0); -- 
    -- CP-element group 28:  transition  input  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Sample/ra
      -- 
    ra_421_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_134_inst_ack_0, ack => testConfigure_CP_0_elements(28)); -- 
    -- CP-element group 29:  transition  input  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	249 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/ca
      -- 
    ca_426_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_134_inst_ack_1, ack => testConfigure_CP_0_elements(29)); -- 
    -- CP-element group 30:  transition  delay-element  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	21 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	23 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_ptr_deref_122_delay
      -- 
    -- Element group testConfigure_CP_0_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(21), ack => testConfigure_CP_0_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  branch  join  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	16 
    -- CP-element group 31: 	17 
    -- CP-element group 31: 	22 
    -- CP-element group 31: 	25 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	32 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (10) 
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135__exit__
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136__entry__
      -- CP-element group 31: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_dead_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/$exit
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_eval_test/branch_req
      -- CP-element group 31: 	 branch_block_stmt_32/R_cmp_137_place
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_if_link/$entry
      -- CP-element group 31: 	 branch_block_stmt_32/if_stmt_136_else_link/$entry
      -- 
    branch_req_435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(31), ack => if_stmt_136_branch_req_0); -- 
    testConfigure_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(16) & testConfigure_CP_0_elements(17) & testConfigure_CP_0_elements(22) & testConfigure_CP_0_elements(25) & testConfigure_CP_0_elements(29);
      gj_testConfigure_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  fork  transition  place  input  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	31 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	234 
    -- CP-element group 32: 	235 
    -- CP-element group 32: 	237 
    -- CP-element group 32: 	238 
    -- CP-element group 32:  members (20) 
      -- CP-element group 32: 	 branch_block_stmt_32/if_stmt_136_if_link/$exit
      -- CP-element group 32: 	 branch_block_stmt_32/if_stmt_136_if_link/if_choice_transition
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/cr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/cr
      -- 
    if_choice_transition_440_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_136_branch_ack_1, ack => testConfigure_CP_0_elements(32)); -- 
    rr_2663_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2663_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_76_inst_req_0); -- 
    cr_2668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_76_inst_req_1); -- 
    rr_2686_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2686_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_83_inst_req_0); -- 
    cr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2691_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(32), ack => type_cast_83_inst_req_1); -- 
    -- CP-element group 33:  fork  transition  place  input  output  bypass 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	250 
    -- CP-element group 33: 	251 
    -- CP-element group 33:  members (12) 
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_136_else_link/$exit
      -- CP-element group 33: 	 branch_block_stmt_32/if_stmt_136_else_link/else_choice_transition
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/rr
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/cr
      -- 
    else_choice_transition_444_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_136_branch_ack_0, ack => testConfigure_CP_0_elements(33)); -- 
    rr_2756_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2756_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_146_inst_req_0); -- 
    cr_2761_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2761_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(33), ack => type_cast_146_inst_req_1); -- 
    -- CP-element group 34:  transition  input  bypass 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	261 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (5) 
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/$exit
      -- CP-element group 34: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/ra
      -- 
    ra_488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_164_store_0_ack_0, ack => testConfigure_CP_0_elements(34)); -- 
    -- CP-element group 35:  branch  transition  place  input  output  bypass 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	261 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	36 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (15) 
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172__exit__
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173__entry__
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/ca
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_dead_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/$exit
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_eval_test/branch_req
      -- CP-element group 35: 	 branch_block_stmt_32/R_cmp12223_174_place
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_if_link/$entry
      -- CP-element group 35: 	 branch_block_stmt_32/if_stmt_173_else_link/$entry
      -- 
    ca_499_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_164_store_0_ack_1, ack => testConfigure_CP_0_elements(35)); -- 
    branch_req_507_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_507_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(35), ack => if_stmt_173_branch_req_0); -- 
    -- CP-element group 36:  transition  place  input  bypass 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	35 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	268 
    -- CP-element group 36:  members (5) 
      -- CP-element group 36: 	 branch_block_stmt_32/if_stmt_173_if_link/$exit
      -- CP-element group 36: 	 branch_block_stmt_32/if_stmt_173_if_link/if_choice_transition
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph221
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph221_PhiReq/$entry
      -- CP-element group 36: 	 branch_block_stmt_32/forx_xend_bbx_xnph221_PhiReq/$exit
      -- 
    if_choice_transition_512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_173_branch_ack_1, ack => testConfigure_CP_0_elements(36)); -- 
    -- CP-element group 37:  merge  transition  place  input  bypass 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	265 
    -- CP-element group 37:  members (14) 
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179__exit__
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_173_else_link/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/if_stmt_173_else_link/else_choice_transition
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xend_forx_xbody14x_xpreheader_PhiReq/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiReqMerge
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/$exit
      -- CP-element group 37: 	 branch_block_stmt_32/merge_stmt_179_PhiAck/dummy
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/$entry
      -- CP-element group 37: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$entry
      -- 
    else_choice_transition_516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_173_branch_ack_0, ack => testConfigure_CP_0_elements(37)); -- 
    -- CP-element group 38:  transition  input  bypass 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	267 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/ra
      -- 
    ra_530_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_198_inst_ack_0, ack => testConfigure_CP_0_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	267 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	55 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_update_completed_
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/ca
      -- 
    ca_535_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_198_inst_ack_1, ack => testConfigure_CP_0_elements(39)); -- 
    -- CP-element group 40:  transition  input  bypass 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	267 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	55 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_sample_complete
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/ack
      -- 
    ack_561_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_204_index_offset_ack_0, ack => testConfigure_CP_0_elements(40)); -- 
    -- CP-element group 41:  transition  input  output  bypass 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	267 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	42 
    -- CP-element group 41:  members (11) 
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_root_address_calculated
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_offset_calculated
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/ack
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/$exit
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/sum_rename_req
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_base_plus_offset/sum_rename_ack
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/$entry
      -- CP-element group 41: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/req
      -- 
    ack_566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_204_index_offset_ack_1, ack => testConfigure_CP_0_elements(41)); -- 
    req_575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(41), ack => addr_of_205_final_reg_req_0); -- 
    -- CP-element group 42:  transition  input  bypass 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/$exit
      -- CP-element group 42: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_request/ack
      -- 
    ack_576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_205_final_reg_ack_0, ack => testConfigure_CP_0_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	267 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	48 
    -- CP-element group 43:  members (19) 
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_root_address_calculated
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_address_resized
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/base_resize_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_addr_resize/base_resize_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/sum_rename_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_base_plus_offset/sum_rename_ack
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/$entry
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/$exit
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/root_register_req
      -- CP-element group 43: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_word_addrgen/root_register_ack
      -- 
    ack_581_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_205_final_reg_ack_1, ack => testConfigure_CP_0_elements(43)); -- 
    -- CP-element group 44:  transition  input  output  bypass 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	267 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	45 
    -- CP-element group 44:  members (6) 
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_update_start_
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/ra
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/$entry
      -- CP-element group 44: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/cr
      -- 
    ra_590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_208_inst_ack_0, ack => testConfigure_CP_0_elements(44)); -- 
    cr_594_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_594_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(44), ack => RPIPE_ConvTranspose_input_pipe_208_inst_req_1); -- 
    -- CP-element group 45:  transition  input  output  bypass 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	44 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	46 
    -- CP-element group 45:  members (6) 
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Update/ca
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/rr
      -- 
    ca_595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_208_inst_ack_1, ack => testConfigure_CP_0_elements(45)); -- 
    rr_603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(45), ack => type_cast_212_inst_req_0); -- 
    -- CP-element group 46:  transition  input  bypass 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/$exit
      -- CP-element group 46: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Sample/ra
      -- 
    ra_604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_0, ack => testConfigure_CP_0_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	267 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_update_completed_
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/ca
      -- 
    ca_609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_212_inst_ack_1, ack => testConfigure_CP_0_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	47 
    -- CP-element group 48: 	43 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48:  members (9) 
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/$exit
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/split_req
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/ptr_deref_215_Split/split_ack
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/$entry
      -- CP-element group 48: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/rr
      -- 
    rr_647_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_647_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(48), ack => ptr_deref_215_store_0_req_0); -- 
    testConfigure_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(47) & testConfigure_CP_0_elements(43);
      gj_testConfigure_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  transition  input  bypass 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	48 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	54 
    -- CP-element group 49:  members (5) 
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/$exit
      -- CP-element group 49: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Sample/word_access_start/word_0/ra
      -- 
    ra_648_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_215_store_0_ack_0, ack => testConfigure_CP_0_elements(49)); -- 
    -- CP-element group 50:  transition  input  bypass 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	267 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	55 
    -- CP-element group 50:  members (5) 
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_update_completed_
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/$exit
      -- CP-element group 50: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/ca
      -- 
    ca_659_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_215_store_0_ack_1, ack => testConfigure_CP_0_elements(50)); -- 
    -- CP-element group 51:  join  transition  output  bypass 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	54 
    -- CP-element group 51: 	267 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	52 
    -- CP-element group 51:  members (5) 
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/$entry
      -- CP-element group 51: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/rr
      -- 
    rr_692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(51), ack => ptr_deref_232_load_0_req_0); -- 
    testConfigure_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(54) & testConfigure_CP_0_elements(267);
      gj_testConfigure_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  transition  input  bypass 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	51 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (5) 
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/$exit
      -- CP-element group 52: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Sample/word_access_start/word_0/ra
      -- 
    ra_693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_232_load_0_ack_0, ack => testConfigure_CP_0_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	267 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (9) 
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/ca
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/$entry
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/$exit
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/merge_req
      -- CP-element group 53: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/ptr_deref_232_Merge/merge_ack
      -- 
    ca_704_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_232_load_0_ack_1, ack => testConfigure_CP_0_elements(53)); -- 
    -- CP-element group 54:  transition  delay-element  bypass 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	49 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	51 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_ptr_deref_232_delay
      -- 
    -- Element group testConfigure_CP_0_elements(54) is a control-delay.
    cp_element_54_delay: control_delay_element  generic map(name => " 54_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(49), ack => testConfigure_CP_0_elements(54), clk => clk, reset =>reset);
    -- CP-element group 55:  branch  join  transition  place  output  bypass 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	40 
    -- CP-element group 55: 	39 
    -- CP-element group 55: 	50 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (10) 
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238__exit__
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239__entry__
      -- CP-element group 55: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_dead_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/$exit
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_eval_test/branch_req
      -- CP-element group 55: 	 branch_block_stmt_32/R_cmp12_240_place
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_if_link/$entry
      -- CP-element group 55: 	 branch_block_stmt_32/if_stmt_239_else_link/$entry
      -- 
    branch_req_718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(55), ack => if_stmt_239_branch_req_0); -- 
    testConfigure_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(40) & testConfigure_CP_0_elements(39) & testConfigure_CP_0_elements(50) & testConfigure_CP_0_elements(53);
      gj_testConfigure_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  place  input  output  bypass 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	262 
    -- CP-element group 56: 	263 
    -- CP-element group 56:  members (12) 
      -- CP-element group 56: 	 branch_block_stmt_32/if_stmt_239_if_link/$exit
      -- CP-element group 56: 	 branch_block_stmt_32/if_stmt_239_if_link/if_choice_transition
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/rr
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/$entry
      -- CP-element group 56: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/cr
      -- 
    if_choice_transition_723_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_239_branch_ack_1, ack => testConfigure_CP_0_elements(56)); -- 
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2856_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_185_inst_req_0); -- 
    cr_2861_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2861_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(56), ack => type_cast_185_inst_req_1); -- 
    -- CP-element group 57:  merge  transition  place  input  bypass 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	268 
    -- CP-element group 57:  members (13) 
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245__exit__
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph221x_xloopexit_bbx_xnph221
      -- CP-element group 57: 	 branch_block_stmt_32/if_stmt_239_else_link/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/if_stmt_239_else_link/else_choice_transition
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph221x_xloopexit
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/forx_xbody14_bbx_xnph221x_xloopexit_PhiReq/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiReqMerge
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/$exit
      -- CP-element group 57: 	 branch_block_stmt_32/merge_stmt_245_PhiAck/dummy
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$entry
      -- CP-element group 57: 	 branch_block_stmt_32/bbx_xnph221x_xloopexit_bbx_xnph221_PhiReq/$exit
      -- 
    else_choice_transition_727_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_239_branch_ack_0, ack => testConfigure_CP_0_elements(57)); -- 
    -- CP-element group 58:  transition  input  output  bypass 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	268 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_update_start_
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/ra
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/cr
      -- 
    ra_741_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_249_inst_ack_0, ack => testConfigure_CP_0_elements(58)); -- 
    cr_745_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_745_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(58), ack => RPIPE_ConvTranspose_input_pipe_249_inst_req_1); -- 
    -- CP-element group 59:  transition  input  output  bypass 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	60 
    -- CP-element group 59:  members (6) 
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Update/ca
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/rr
      -- 
    ca_746_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_249_inst_ack_1, ack => testConfigure_CP_0_elements(59)); -- 
    rr_754_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_754_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(59), ack => type_cast_253_inst_req_0); -- 
    -- CP-element group 60:  transition  input  bypass 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	59 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Sample/ra
      -- 
    ra_755_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_0, ack => testConfigure_CP_0_elements(60)); -- 
    -- CP-element group 61:  fork  transition  place  input  output  bypass 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	268 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	269 
    -- CP-element group 61: 	270 
    -- CP-element group 61: 	271 
    -- CP-element group 61:  members (17) 
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254__exit__
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/ca
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/$entry
      -- CP-element group 61: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/cr
      -- 
    ca_760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_253_inst_ack_1, ack => testConfigure_CP_0_elements(61)); -- 
    rr_2929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_267_inst_req_0); -- 
    cr_2934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(61), ack => type_cast_267_inst_req_1); -- 
    -- CP-element group 62:  transition  input  bypass 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	284 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/ack
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/$exit
      -- 
    ack_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_274_final_reg_ack_0, ack => testConfigure_CP_0_elements(62)); -- 
    -- CP-element group 63:  join  fork  transition  input  output  bypass 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	284 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (28) 
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_root_address_calculated
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_address_resized
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/base_resize_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_addr_resize/base_resize_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/sum_rename_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_base_plus_offset/sum_rename_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/root_register_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_word_addrgen/root_register_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/$exit
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/split_req
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/ptr_deref_277_Split/split_ack
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/$entry
      -- CP-element group 63: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/rr
      -- 
    ack_802_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_274_final_reg_ack_1, ack => testConfigure_CP_0_elements(63)); -- 
    rr_840_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_840_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(63), ack => ptr_deref_277_store_0_req_0); -- 
    -- CP-element group 64:  transition  input  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	63 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (5) 
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/$exit
      -- CP-element group 64: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Sample/word_access_start/word_0/ra
      -- 
    ra_841_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_277_store_0_ack_0, ack => testConfigure_CP_0_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	284 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	70 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/$exit
      -- CP-element group 65: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/ca
      -- 
    ca_852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_277_store_0_ack_1, ack => testConfigure_CP_0_elements(65)); -- 
    -- CP-element group 66:  transition  input  output  bypass 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	284 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_update_start_
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/ra
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/cr
      -- 
    ra_861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_0, ack => testConfigure_CP_0_elements(66)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(66), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_1); -- 
    -- CP-element group 67:  transition  input  output  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (6) 
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Update/ca
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/rr
      -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_281_inst_ack_1, ack => testConfigure_CP_0_elements(67)); -- 
    rr_874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(67), ack => type_cast_285_inst_req_0); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Sample/ra
      -- 
    ra_875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_0, ack => testConfigure_CP_0_elements(68)); -- 
    -- CP-element group 69:  transition  input  bypass 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	284 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	70 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/ca
      -- 
    ca_880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_285_inst_ack_1, ack => testConfigure_CP_0_elements(69)); -- 
    -- CP-element group 70:  branch  join  transition  place  output  bypass 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	65 
    -- CP-element group 70: 	69 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (10) 
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298__exit__
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299__entry__
      -- CP-element group 70: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_dead_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/$exit
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_eval_test/branch_req
      -- CP-element group 70: 	 branch_block_stmt_32/R_exitcond_300_place
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_if_link/$entry
      -- CP-element group 70: 	 branch_block_stmt_32/if_stmt_299_else_link/$entry
      -- 
    branch_req_888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(70), ack => if_stmt_299_branch_req_0); -- 
    testConfigure_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(65) & testConfigure_CP_0_elements(69);
      gj_testConfigure_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  place  input  output  bypass 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	285 
    -- CP-element group 71: 	286 
    -- CP-element group 71:  members (12) 
      -- CP-element group 71: 	 branch_block_stmt_32/if_stmt_299_if_link/$exit
      -- CP-element group 71: 	 branch_block_stmt_32/if_stmt_299_if_link/if_choice_transition
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/rr
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/cr
      -- 
    if_choice_transition_893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_1, ack => testConfigure_CP_0_elements(71)); -- 
    rr_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_309_inst_req_0); -- 
    cr_3019_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3019_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(71), ack => type_cast_309_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  place  input  output  bypass 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	274 
    -- CP-element group 72: 	275 
    -- CP-element group 72: 	277 
    -- CP-element group 72: 	278 
    -- CP-element group 72:  members (20) 
      -- CP-element group 72: 	 branch_block_stmt_32/if_stmt_299_else_link/$exit
      -- CP-element group 72: 	 branch_block_stmt_32/if_stmt_299_else_link/else_choice_transition
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/cr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/rr
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/$entry
      -- CP-element group 72: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/cr
      -- 
    else_choice_transition_897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_299_branch_ack_0, ack => testConfigure_CP_0_elements(72)); -- 
    rr_2955_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2955_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_263_inst_req_0); -- 
    cr_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_263_inst_req_1); -- 
    rr_2978_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2978_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_269_inst_req_0); -- 
    cr_2983_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2983_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(72), ack => type_cast_269_inst_req_1); -- 
    -- CP-element group 73:  join  fork  transition  output  bypass 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	288 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73: 	75 
    -- CP-element group 73: 	76 
    -- CP-element group 73: 	79 
    -- CP-element group 73: 	80 
    -- CP-element group 73: 	82 
    -- CP-element group 73: 	86 
    -- CP-element group 73: 	87 
    -- CP-element group 73: 	89 
    -- CP-element group 73: 	93 
    -- CP-element group 73: 	94 
    -- CP-element group 73: 	96 
    -- CP-element group 73: 	97 
    -- CP-element group 73: 	98 
    -- CP-element group 73: 	99 
    -- CP-element group 73: 	100 
    -- CP-element group 73: 	101 
    -- CP-element group 73: 	102 
    -- CP-element group 73: 	105 
    -- CP-element group 73: 	106 
    -- CP-element group 73: 	107 
    -- CP-element group 73: 	108 
    -- CP-element group 73: 	109 
    -- CP-element group 73: 	110 
    -- CP-element group 73: 	111 
    -- CP-element group 73: 	112 
    -- CP-element group 73: 	113 
    -- CP-element group 73: 	116 
    -- CP-element group 73:  members (280) 
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/split_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/STORE_padding_311_Split/split_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/rr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/cr
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_update_start_
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_root_address_calculated
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_address_resized
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/base_resize_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_addr_resize/base_resize_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/sum_rename_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_base_plus_offset/sum_rename_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/$exit
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/root_register_req
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_word_addrgen/root_register_ack
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/$entry
      -- CP-element group 73: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/cr
      -- 
    cr_934_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_934_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_311_store_0_req_1); -- 
    rr_923_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_923_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => STORE_padding_311_store_0_req_0); -- 
    rr_943_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_943_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => RPIPE_ConvTranspose_input_pipe_315_inst_req_0); -- 
    cr_962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_319_inst_req_1); -- 
    cr_1012_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1012_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_330_store_0_req_1); -- 
    cr_1040_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1040_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_338_inst_req_1); -- 
    cr_1090_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1090_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_349_store_0_req_1); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1118_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_357_inst_req_1); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_368_store_0_req_1); -- 
    cr_1213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_381_load_0_req_1); -- 
    rr_1202_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1202_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_381_load_0_req_0); -- 
    cr_1263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_393_load_0_req_1); -- 
    rr_1252_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1252_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_393_load_0_req_0); -- 
    cr_1313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_405_load_0_req_1); -- 
    rr_1302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_405_load_0_req_0); -- 
    cr_1332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_419_inst_req_1); -- 
    cr_1377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_431_load_0_req_1); -- 
    rr_1366_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1366_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_431_load_0_req_0); -- 
    cr_1427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_443_load_0_req_1); -- 
    rr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_443_load_0_req_0); -- 
    cr_1477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_455_load_0_req_1); -- 
    rr_1466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_455_load_0_req_0); -- 
    cr_1527_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1527_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_467_load_0_req_1); -- 
    rr_1516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => ptr_deref_467_load_0_req_0); -- 
    cr_1546_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1546_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(73), ack => type_cast_486_inst_req_1); -- 
    testConfigure_CP_0_elements(73) <= testConfigure_CP_0_elements(288);
    -- CP-element group 74:  transition  input  bypass 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (5) 
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/$exit
      -- CP-element group 74: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Sample/word_access_start/word_0/ra
      -- 
    ra_924_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_311_store_0_ack_0, ack => testConfigure_CP_0_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	119 
    -- CP-element group 75:  members (5) 
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/$exit
      -- CP-element group 75: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/STORE_padding_311_Update/word_access_complete/word_0/ca
      -- 
    ca_935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => STORE_padding_311_store_0_ack_1, ack => testConfigure_CP_0_elements(75)); -- 
    -- CP-element group 76:  transition  input  output  bypass 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	73 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	77 
    -- CP-element group 76:  members (6) 
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_update_start_
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Sample/ra
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/$entry
      -- CP-element group 76: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/cr
      -- 
    ra_944_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_315_inst_ack_0, ack => testConfigure_CP_0_elements(76)); -- 
    cr_948_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_948_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(76), ack => RPIPE_ConvTranspose_input_pipe_315_inst_req_1); -- 
    -- CP-element group 77:  fork  transition  input  output  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	76 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77: 	83 
    -- CP-element group 77:  members (9) 
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_315_Update/ca
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/rr
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/rr
      -- 
    ca_949_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_315_inst_ack_1, ack => testConfigure_CP_0_elements(77)); -- 
    rr_957_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_957_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => type_cast_319_inst_req_0); -- 
    rr_1021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(77), ack => RPIPE_ConvTranspose_input_pipe_334_inst_req_0); -- 
    -- CP-element group 78:  transition  input  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Sample/ra
      -- 
    ra_958_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_0, ack => testConfigure_CP_0_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	73 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_319_Update/ca
      -- 
    ca_963_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_319_inst_ack_1, ack => testConfigure_CP_0_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	73 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (9) 
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/$exit
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/split_req
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/ptr_deref_330_Split/split_ack
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/$entry
      -- CP-element group 80: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/rr
      -- 
    rr_1001_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1001_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(80), ack => ptr_deref_330_store_0_req_0); -- 
    testConfigure_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(79);
      gj_testConfigure_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  transition  input  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	117 
    -- CP-element group 81:  members (5) 
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/$exit
      -- CP-element group 81: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Sample/word_access_start/word_0/ra
      -- 
    ra_1002_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_330_store_0_ack_0, ack => testConfigure_CP_0_elements(81)); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	73 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	119 
    -- CP-element group 82:  members (5) 
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/$exit
      -- CP-element group 82: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_Update/word_access_complete/word_0/ca
      -- 
    ca_1013_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_330_store_0_ack_1, ack => testConfigure_CP_0_elements(82)); -- 
    -- CP-element group 83:  transition  input  output  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	77 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	84 
    -- CP-element group 83:  members (6) 
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_update_start_
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/$exit
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/cr
      -- 
    ra_1022_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_334_inst_ack_0, ack => testConfigure_CP_0_elements(83)); -- 
    cr_1026_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1026_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(83), ack => RPIPE_ConvTranspose_input_pipe_334_inst_req_1); -- 
    -- CP-element group 84:  fork  transition  input  output  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	83 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84: 	90 
    -- CP-element group 84:  members (9) 
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_334_Update/ca
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/rr
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/rr
      -- 
    ca_1027_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_334_inst_ack_1, ack => testConfigure_CP_0_elements(84)); -- 
    rr_1035_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1035_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => type_cast_338_inst_req_0); -- 
    rr_1099_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1099_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(84), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_0); -- 
    -- CP-element group 85:  transition  input  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Sample/ra
      -- 
    ra_1036_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_0, ack => testConfigure_CP_0_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	73 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_338_Update/ca
      -- 
    ca_1041_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_1, ack => testConfigure_CP_0_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	73 
    -- CP-element group 87: 	86 
    -- CP-element group 87: 	117 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (9) 
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/$exit
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/split_req
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/ptr_deref_349_Split/split_ack
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/$entry
      -- CP-element group 87: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/rr
      -- 
    rr_1079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(87), ack => ptr_deref_349_store_0_req_0); -- 
    testConfigure_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(86) & testConfigure_CP_0_elements(117);
      gj_testConfigure_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	87 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	118 
    -- CP-element group 88:  members (5) 
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_sample_completed_
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/$exit
      -- CP-element group 88: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Sample/word_access_start/word_0/ra
      -- 
    ra_1080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_store_0_ack_0, ack => testConfigure_CP_0_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	73 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	119 
    -- CP-element group 89:  members (5) 
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_update_completed_
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/$exit
      -- CP-element group 89: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_Update/word_access_complete/word_0/ca
      -- 
    ca_1091_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_349_store_0_ack_1, ack => testConfigure_CP_0_elements(89)); -- 
    -- CP-element group 90:  transition  input  output  bypass 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	84 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	91 
    -- CP-element group 90:  members (6) 
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_update_start_
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Sample/ra
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/$entry
      -- CP-element group 90: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/cr
      -- 
    ra_1100_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_0, ack => testConfigure_CP_0_elements(90)); -- 
    cr_1104_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1104_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(90), ack => RPIPE_ConvTranspose_input_pipe_353_inst_req_1); -- 
    -- CP-element group 91:  transition  input  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	90 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	92 
    -- CP-element group 91:  members (6) 
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/RPIPE_ConvTranspose_input_pipe_353_Update/ca
      -- CP-element group 91: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_sample_start_
      -- 
    ca_1105_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_353_inst_ack_1, ack => testConfigure_CP_0_elements(91)); -- 
    rr_1113_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1113_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(91), ack => type_cast_357_inst_req_0); -- 
    -- CP-element group 92:  transition  input  bypass 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	91 
    -- CP-element group 92: successors 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/ra
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_sample_completed_
      -- 
    ra_1114_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_0, ack => testConfigure_CP_0_elements(92)); -- 
    -- CP-element group 93:  transition  input  bypass 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	73 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	94 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/ca
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_357_update_completed_
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_357_inst_ack_1, ack => testConfigure_CP_0_elements(93)); -- 
    -- CP-element group 94:  join  transition  output  bypass 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	73 
    -- CP-element group 94: 	93 
    -- CP-element group 94: 	118 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	95 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_sample_start_
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/rr
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/split_ack
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/split_req
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/$exit
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/ptr_deref_368_Split/$entry
      -- CP-element group 94: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/$entry
      -- 
    rr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(94), ack => ptr_deref_368_store_0_req_0); -- 
    testConfigure_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "testConfigure_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(73) & testConfigure_CP_0_elements(93) & testConfigure_CP_0_elements(118);
      gj_testConfigure_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  transition  input  bypass 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	94 
    -- CP-element group 95: successors 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_sample_completed_
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/ra
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/word_0/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/word_access_start/$exit
      -- CP-element group 95: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Sample/$exit
      -- 
    ra_1158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_368_store_0_ack_0, ack => testConfigure_CP_0_elements(95)); -- 
    -- CP-element group 96:  transition  input  bypass 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	73 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	119 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/ca
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/word_0/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/word_access_complete/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_Update/$exit
      -- CP-element group 96: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_368_update_completed_
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 96_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_368_store_0_ack_1, ack => testConfigure_CP_0_elements(96)); -- 
    -- CP-element group 97:  transition  input  bypass 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	73 
    -- CP-element group 97: successors 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/word_0/ra
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Sample/$exit
      -- 
    ra_1203_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_load_0_ack_0, ack => testConfigure_CP_0_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	73 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	103 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/merge_ack
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/ptr_deref_381_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/word_access_complete/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_381_update_completed_
      -- 
    ca_1214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_381_load_0_ack_1, ack => testConfigure_CP_0_elements(98)); -- 
    -- CP-element group 99:  transition  input  bypass 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	73 
    -- CP-element group 99: successors 
    -- CP-element group 99:  members (5) 
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/$exit
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_sample_completed_
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/ra
      -- CP-element group 99: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Sample/word_access_start/word_0/$exit
      -- 
    ra_1253_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_393_load_0_ack_0, ack => testConfigure_CP_0_elements(99)); -- 
    -- CP-element group 100:  transition  input  bypass 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	73 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	103 
    -- CP-element group 100:  members (9) 
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/merge_ack
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/merge_req
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/ptr_deref_393_Merge/$entry
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/ca
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/word_0/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_update_completed_
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/word_access_complete/$exit
      -- CP-element group 100: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_393_Update/$exit
      -- 
    ca_1264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_393_load_0_ack_1, ack => testConfigure_CP_0_elements(100)); -- 
    -- CP-element group 101:  transition  input  bypass 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	73 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (5) 
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/ra
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/word_0/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/word_access_start/$exit
      -- CP-element group 101: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Sample/$exit
      -- 
    ra_1303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_0, ack => testConfigure_CP_0_elements(101)); -- 
    -- CP-element group 102:  transition  input  bypass 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	73 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	103 
    -- CP-element group 102:  members (9) 
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/merge_ack
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/merge_req
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/ptr_deref_405_Merge/$entry
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/ca
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/word_0/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/word_access_complete/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_405_update_completed_
      -- 
    ca_1314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_405_load_0_ack_1, ack => testConfigure_CP_0_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	98 
    -- CP-element group 103: 	100 
    -- CP-element group 103: 	102 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	104 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/rr
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_sample_start_
      -- 
    rr_1327_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1327_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(103), ack => type_cast_419_inst_req_0); -- 
    testConfigure_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(98) & testConfigure_CP_0_elements(100) & testConfigure_CP_0_elements(102);
      gj_testConfigure_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  transition  input  bypass 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	103 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/ra
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_sample_completed_
      -- 
    ra_1328_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_0, ack => testConfigure_CP_0_elements(104)); -- 
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	73 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	119 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/ca
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_419_update_completed_
      -- 
    ca_1333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_419_inst_ack_1, ack => testConfigure_CP_0_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	73 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_sample_completed_
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/ra
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/word_0/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/word_access_start/$exit
      -- CP-element group 106: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Sample/$exit
      -- 
    ra_1367_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_load_0_ack_0, ack => testConfigure_CP_0_elements(106)); -- 
    -- CP-element group 107:  transition  input  bypass 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	73 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	114 
    -- CP-element group 107:  members (9) 
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/merge_ack
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_update_completed_
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/merge_req
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/$exit
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/ptr_deref_431_Merge/$entry
      -- CP-element group 107: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_431_Update/word_access_complete/word_0/ca
      -- 
    ca_1378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 107_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_431_load_0_ack_1, ack => testConfigure_CP_0_elements(107)); -- 
    -- CP-element group 108:  transition  input  bypass 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	73 
    -- CP-element group 108: successors 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_sample_completed_
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/ra
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/word_0/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/word_access_start/$exit
      -- CP-element group 108: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Sample/$exit
      -- 
    ra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 108_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_443_load_0_ack_0, ack => testConfigure_CP_0_elements(108)); -- 
    -- CP-element group 109:  transition  input  bypass 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	73 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	114 
    -- CP-element group 109:  members (9) 
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/merge_ack
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/merge_req
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/ptr_deref_443_Merge/$entry
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/ca
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/word_0/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/word_access_complete/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_Update/$exit
      -- CP-element group 109: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_443_update_completed_
      -- 
    ca_1428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_443_load_0_ack_1, ack => testConfigure_CP_0_elements(109)); -- 
    -- CP-element group 110:  transition  input  bypass 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	73 
    -- CP-element group 110: successors 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/ra
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Sample/$exit
      -- 
    ra_1467_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_455_load_0_ack_0, ack => testConfigure_CP_0_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	73 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	114 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/merge_ack
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/ptr_deref_455_Merge/$entry
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_455_Update/$exit
      -- 
    ca_1478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_455_load_0_ack_1, ack => testConfigure_CP_0_elements(111)); -- 
    -- CP-element group 112:  transition  input  bypass 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	73 
    -- CP-element group 112: successors 
    -- CP-element group 112:  members (5) 
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/ra
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/word_0/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Sample/word_access_start/$exit
      -- 
    ra_1517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_0, ack => testConfigure_CP_0_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	73 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (9) 
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/$entry
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/ca
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/merge_ack
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/word_0/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/ptr_deref_467_Merge/merge_req
      -- CP-element group 113: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_467_Update/word_access_complete/$exit
      -- 
    ca_1528_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_1, ack => testConfigure_CP_0_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	107 
    -- CP-element group 114: 	109 
    -- CP-element group 114: 	111 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/rr
      -- CP-element group 114: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/$entry
      -- 
    rr_1541_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1541_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(114), ack => type_cast_486_inst_req_0); -- 
    testConfigure_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(107) & testConfigure_CP_0_elements(109) & testConfigure_CP_0_elements(111) & testConfigure_CP_0_elements(113);
      gj_testConfigure_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  transition  input  bypass 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/ra
      -- CP-element group 115: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Sample/$exit
      -- 
    ra_1542_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_0, ack => testConfigure_CP_0_elements(115)); -- 
    -- CP-element group 116:  transition  input  bypass 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	73 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	119 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/ca
      -- CP-element group 116: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/type_cast_486_Update/$exit
      -- 
    ca_1547_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_486_inst_ack_1, ack => testConfigure_CP_0_elements(116)); -- 
    -- CP-element group 117:  transition  delay-element  bypass 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	81 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	87 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_330_ptr_deref_349_delay
      -- 
    -- Element group testConfigure_CP_0_elements(117) is a control-delay.
    cp_element_117_delay: control_delay_element  generic map(name => " 117_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(81), ack => testConfigure_CP_0_elements(117), clk => clk, reset =>reset);
    -- CP-element group 118:  transition  delay-element  bypass 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	88 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	94 
    -- CP-element group 118:  members (1) 
      -- CP-element group 118: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/ptr_deref_349_ptr_deref_368_delay
      -- 
    -- Element group testConfigure_CP_0_elements(118) is a control-delay.
    cp_element_118_delay: control_delay_element  generic map(name => " 118_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(88), ack => testConfigure_CP_0_elements(118), clk => clk, reset =>reset);
    -- CP-element group 119:  branch  join  transition  place  output  bypass 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	75 
    -- CP-element group 119: 	82 
    -- CP-element group 119: 	89 
    -- CP-element group 119: 	96 
    -- CP-element group 119: 	105 
    -- CP-element group 119: 	116 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	120 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (10) 
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_dead_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/R_cmp65213_501_place
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_if_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_else_link/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/$entry
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/$exit
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500_eval_test/branch_req
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499__exit__
      -- CP-element group 119: 	 branch_block_stmt_32/if_stmt_500__entry__
      -- CP-element group 119: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499/$exit
      -- 
    branch_req_1557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(119), ack => if_stmt_500_branch_req_0); -- 
    testConfigure_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(75) & testConfigure_CP_0_elements(82) & testConfigure_CP_0_elements(89) & testConfigure_CP_0_elements(96) & testConfigure_CP_0_elements(105) & testConfigure_CP_0_elements(116);
      gj_testConfigure_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  transition  place  input  bypass 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	119 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	289 
    -- CP-element group 120:  members (5) 
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_500_if_link/$exit
      -- CP-element group 120: 	 branch_block_stmt_32/if_stmt_500_if_link/if_choice_transition
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 120: 	 branch_block_stmt_32/forx_xend37_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_1, ack => testConfigure_CP_0_elements(120)); -- 
    -- CP-element group 121:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	124 
    -- CP-element group 121: 	125 
    -- CP-element group 121:  members (18) 
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_500_else_link/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/if_stmt_500_else_link/else_choice_transition
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph215
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527__exit__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560__entry__
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_update_start_
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/rr
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/cr
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph215_PhiReq/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/forx_xend37_bbx_xnph215_PhiReq/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiReqMerge
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/$entry
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/$exit
      -- CP-element group 121: 	 branch_block_stmt_32/merge_stmt_527_PhiAck/dummy
      -- 
    else_choice_transition_1566_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_500_branch_ack_0, ack => testConfigure_CP_0_elements(121)); -- 
    rr_1601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_540_inst_req_0); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1606_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(121), ack => type_cast_540_inst_req_1); -- 
    -- CP-element group 122:  transition  place  input  bypass 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	289 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	302 
    -- CP-element group 122:  members (5) 
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_521_if_link/$exit
      -- CP-element group 122: 	 branch_block_stmt_32/if_stmt_521_if_link/if_choice_transition
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$entry
      -- CP-element group 122: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_1584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_521_branch_ack_1, ack => testConfigure_CP_0_elements(122)); -- 
    -- CP-element group 123:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	289 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	168 
    -- CP-element group 123: 	169 
    -- CP-element group 123:  members (18) 
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732__exit__
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770__entry__
      -- CP-element group 123: 	 branch_block_stmt_32/if_stmt_521_else_link/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/if_stmt_521_else_link/else_choice_transition
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph210
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_update_start_
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/rr
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/cr
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/forx_xcond119x_xpreheader_bbx_xnph210_PhiReq/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiReqMerge
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/$entry
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/$exit
      -- CP-element group 123: 	 branch_block_stmt_32/merge_stmt_732_PhiAck/dummy
      -- 
    else_choice_transition_1588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_521_branch_ack_0, ack => testConfigure_CP_0_elements(123)); -- 
    rr_1960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_750_inst_req_0); -- 
    cr_1965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(123), ack => type_cast_750_inst_req_1); -- 
    -- CP-element group 124:  transition  input  bypass 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	121 
    -- CP-element group 124: successors 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_sample_completed_
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/$exit
      -- CP-element group 124: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Sample/ra
      -- 
    ra_1602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_0, ack => testConfigure_CP_0_elements(124)); -- 
    -- CP-element group 125:  transition  place  input  bypass 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	121 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	290 
    -- CP-element group 125:  members (9) 
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560__exit__
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_update_completed_
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/$exit
      -- CP-element group 125: 	 branch_block_stmt_32/assign_stmt_532_to_assign_stmt_560/type_cast_540_Update/ca
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/$entry
      -- CP-element group 125: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$entry
      -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_540_inst_ack_1, ack => testConfigure_CP_0_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	295 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	165 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_sample_complete
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/$exit
      -- CP-element group 126: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/ack
      -- 
    ack_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_575_index_offset_ack_0, ack => testConfigure_CP_0_elements(126)); -- 
    -- CP-element group 127:  transition  input  output  bypass 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	295 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	128 
    -- CP-element group 127:  members (11) 
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_root_address_calculated
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_offset_calculated
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/ack
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/$entry
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/$exit
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/sum_rename_req
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_base_plus_offset/sum_rename_ack
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/$entry
      -- CP-element group 127: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/req
      -- 
    ack_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_575_index_offset_ack_1, ack => testConfigure_CP_0_elements(127)); -- 
    req_1650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(127), ack => addr_of_576_final_reg_req_0); -- 
    -- CP-element group 128:  transition  input  bypass 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	127 
    -- CP-element group 128: successors 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_sample_completed_
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/$exit
      -- CP-element group 128: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_request/ack
      -- 
    ack_1651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_576_final_reg_ack_0, ack => testConfigure_CP_0_elements(128)); -- 
    -- CP-element group 129:  fork  transition  input  bypass 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	295 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	162 
    -- CP-element group 129:  members (19) 
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_update_completed_
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_root_address_calculated
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_address_resized
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/base_resize_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_addr_resize/base_resize_ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/sum_rename_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_base_plus_offset/sum_rename_ack
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/$entry
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/$exit
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/root_register_req
      -- CP-element group 129: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_word_addrgen/root_register_ack
      -- 
    ack_1656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_576_final_reg_ack_1, ack => testConfigure_CP_0_elements(129)); -- 
    -- CP-element group 130:  transition  input  output  bypass 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	295 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_update_start_
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/ra
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/cr
      -- 
    ra_1665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_0, ack => testConfigure_CP_0_elements(130)); -- 
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(130), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  output  bypass 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	132 
    -- CP-element group 131: 	134 
    -- CP-element group 131:  members (9) 
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Update/ca
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/rr
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/rr
      -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_579_inst_ack_1, ack => testConfigure_CP_0_elements(131)); -- 
    rr_1678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => type_cast_583_inst_req_0); -- 
    rr_1692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(131), ack => RPIPE_ConvTranspose_input_pipe_592_inst_req_0); -- 
    -- CP-element group 132:  transition  input  bypass 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	131 
    -- CP-element group 132: successors 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_sample_completed_
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/$exit
      -- CP-element group 132: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Sample/ra
      -- 
    ra_1679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 132_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_0, ack => testConfigure_CP_0_elements(132)); -- 
    -- CP-element group 133:  transition  input  bypass 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	295 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	162 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_update_completed_
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/$exit
      -- CP-element group 133: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/ca
      -- 
    ca_1684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_583_inst_ack_1, ack => testConfigure_CP_0_elements(133)); -- 
    -- CP-element group 134:  transition  input  output  bypass 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	131 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	135 
    -- CP-element group 134:  members (6) 
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_update_start_
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Sample/ra
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/$entry
      -- CP-element group 134: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/cr
      -- 
    ra_1693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_592_inst_ack_0, ack => testConfigure_CP_0_elements(134)); -- 
    cr_1697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(134), ack => RPIPE_ConvTranspose_input_pipe_592_inst_req_1); -- 
    -- CP-element group 135:  fork  transition  input  output  bypass 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	134 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135: 	138 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_592_Update/ca
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/rr
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/rr
      -- 
    ca_1698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_592_inst_ack_1, ack => testConfigure_CP_0_elements(135)); -- 
    rr_1706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => type_cast_596_inst_req_0); -- 
    rr_1720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(135), ack => RPIPE_ConvTranspose_input_pipe_610_inst_req_0); -- 
    -- CP-element group 136:  transition  input  bypass 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	135 
    -- CP-element group 136: successors 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_sample_completed_
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/$exit
      -- CP-element group 136: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Sample/ra
      -- 
    ra_1707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 136_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_0, ack => testConfigure_CP_0_elements(136)); -- 
    -- CP-element group 137:  transition  input  bypass 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	295 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	162 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_update_completed_
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/$exit
      -- CP-element group 137: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/ca
      -- 
    ca_1712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_596_inst_ack_1, ack => testConfigure_CP_0_elements(137)); -- 
    -- CP-element group 138:  transition  input  output  bypass 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	135 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	139 
    -- CP-element group 138:  members (6) 
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_sample_completed_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_update_start_
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/$exit
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Sample/ra
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/$entry
      -- CP-element group 138: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/cr
      -- 
    ra_1721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_610_inst_ack_0, ack => testConfigure_CP_0_elements(138)); -- 
    cr_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(138), ack => RPIPE_ConvTranspose_input_pipe_610_inst_req_1); -- 
    -- CP-element group 139:  fork  transition  input  output  bypass 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	138 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	140 
    -- CP-element group 139: 	142 
    -- CP-element group 139:  members (9) 
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_update_completed_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/$exit
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_610_Update/ca
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/rr
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/rr
      -- 
    ca_1726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 139_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_610_inst_ack_1, ack => testConfigure_CP_0_elements(139)); -- 
    rr_1734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => type_cast_614_inst_req_0); -- 
    rr_1748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(139), ack => RPIPE_ConvTranspose_input_pipe_628_inst_req_0); -- 
    -- CP-element group 140:  transition  input  bypass 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	139 
    -- CP-element group 140: successors 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_sample_completed_
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/$exit
      -- CP-element group 140: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Sample/ra
      -- 
    ra_1735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 140_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => testConfigure_CP_0_elements(140)); -- 
    -- CP-element group 141:  transition  input  bypass 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	295 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	162 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_update_completed_
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/$exit
      -- CP-element group 141: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/ca
      -- 
    ca_1740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_1, ack => testConfigure_CP_0_elements(141)); -- 
    -- CP-element group 142:  transition  input  output  bypass 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	143 
    -- CP-element group 142:  members (6) 
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_sample_completed_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_update_start_
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/$exit
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Sample/ra
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/$entry
      -- CP-element group 142: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/cr
      -- 
    ra_1749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_628_inst_ack_0, ack => testConfigure_CP_0_elements(142)); -- 
    cr_1753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(142), ack => RPIPE_ConvTranspose_input_pipe_628_inst_req_1); -- 
    -- CP-element group 143:  fork  transition  input  output  bypass 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	144 
    -- CP-element group 143: 	146 
    -- CP-element group 143:  members (9) 
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_update_completed_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/$exit
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_628_Update/ca
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/rr
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/rr
      -- 
    ca_1754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 143_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_628_inst_ack_1, ack => testConfigure_CP_0_elements(143)); -- 
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => type_cast_632_inst_req_0); -- 
    rr_1776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(143), ack => RPIPE_ConvTranspose_input_pipe_646_inst_req_0); -- 
    -- CP-element group 144:  transition  input  bypass 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: 	143 
    -- CP-element group 144: successors 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_sample_completed_
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/$exit
      -- CP-element group 144: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Sample/ra
      -- 
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 144_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_0, ack => testConfigure_CP_0_elements(144)); -- 
    -- CP-element group 145:  transition  input  bypass 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	295 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	162 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_update_completed_
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/$exit
      -- CP-element group 145: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/ca
      -- 
    ca_1768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_632_inst_ack_1, ack => testConfigure_CP_0_elements(145)); -- 
    -- CP-element group 146:  transition  input  output  bypass 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	143 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	147 
    -- CP-element group 146:  members (6) 
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_sample_completed_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_update_start_
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/$exit
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Sample/ra
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/$entry
      -- CP-element group 146: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/cr
      -- 
    ra_1777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_646_inst_ack_0, ack => testConfigure_CP_0_elements(146)); -- 
    cr_1781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(146), ack => RPIPE_ConvTranspose_input_pipe_646_inst_req_1); -- 
    -- CP-element group 147:  fork  transition  input  output  bypass 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	146 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	148 
    -- CP-element group 147: 	150 
    -- CP-element group 147:  members (9) 
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_update_completed_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/$exit
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_646_Update/ca
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/rr
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/rr
      -- 
    ca_1782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 147_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_646_inst_ack_1, ack => testConfigure_CP_0_elements(147)); -- 
    rr_1790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => type_cast_650_inst_req_0); -- 
    rr_1804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(147), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_0); -- 
    -- CP-element group 148:  transition  input  bypass 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: 	147 
    -- CP-element group 148: successors 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_sample_completed_
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/$exit
      -- CP-element group 148: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Sample/ra
      -- 
    ra_1791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 148_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_0, ack => testConfigure_CP_0_elements(148)); -- 
    -- CP-element group 149:  transition  input  bypass 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	295 
    -- CP-element group 149: successors 
    -- CP-element group 149: 	162 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_update_completed_
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/$exit
      -- CP-element group 149: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/ca
      -- 
    ca_1796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_650_inst_ack_1, ack => testConfigure_CP_0_elements(149)); -- 
    -- CP-element group 150:  transition  input  output  bypass 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	147 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	151 
    -- CP-element group 150:  members (6) 
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_sample_completed_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_update_start_
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/$exit
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Sample/ra
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/$entry
      -- CP-element group 150: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/cr
      -- 
    ra_1805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_0, ack => testConfigure_CP_0_elements(150)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(150), ack => RPIPE_ConvTranspose_input_pipe_664_inst_req_1); -- 
    -- CP-element group 151:  fork  transition  input  output  bypass 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	150 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	152 
    -- CP-element group 151: 	154 
    -- CP-element group 151:  members (9) 
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_update_completed_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/$exit
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_664_Update/ca
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/rr
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/rr
      -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 151_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_664_inst_ack_1, ack => testConfigure_CP_0_elements(151)); -- 
    rr_1818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => type_cast_668_inst_req_0); -- 
    rr_1832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(151), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_0); -- 
    -- CP-element group 152:  transition  input  bypass 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: 	151 
    -- CP-element group 152: successors 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_sample_completed_
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/$exit
      -- CP-element group 152: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Sample/ra
      -- 
    ra_1819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 152_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_0, ack => testConfigure_CP_0_elements(152)); -- 
    -- CP-element group 153:  transition  input  bypass 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	295 
    -- CP-element group 153: successors 
    -- CP-element group 153: 	162 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_update_completed_
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/$exit
      -- CP-element group 153: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/ca
      -- 
    ca_1824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_668_inst_ack_1, ack => testConfigure_CP_0_elements(153)); -- 
    -- CP-element group 154:  transition  input  output  bypass 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	151 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	155 
    -- CP-element group 154:  members (6) 
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_sample_completed_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_update_start_
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/$exit
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Sample/ra
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/$entry
      -- CP-element group 154: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/cr
      -- 
    ra_1833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_0, ack => testConfigure_CP_0_elements(154)); -- 
    cr_1837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(154), ack => RPIPE_ConvTranspose_input_pipe_682_inst_req_1); -- 
    -- CP-element group 155:  fork  transition  input  output  bypass 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	154 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	156 
    -- CP-element group 155: 	158 
    -- CP-element group 155:  members (9) 
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_update_completed_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/$exit
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_682_Update/ca
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/rr
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/rr
      -- 
    ca_1838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 155_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_682_inst_ack_1, ack => testConfigure_CP_0_elements(155)); -- 
    rr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => type_cast_686_inst_req_0); -- 
    rr_1860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(155), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_0); -- 
    -- CP-element group 156:  transition  input  bypass 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: 	155 
    -- CP-element group 156: successors 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_sample_completed_
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/$exit
      -- CP-element group 156: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Sample/ra
      -- 
    ra_1847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 156_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_0, ack => testConfigure_CP_0_elements(156)); -- 
    -- CP-element group 157:  transition  input  bypass 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	295 
    -- CP-element group 157: successors 
    -- CP-element group 157: 	162 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_update_completed_
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/$exit
      -- CP-element group 157: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/ca
      -- 
    ca_1852_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_686_inst_ack_1, ack => testConfigure_CP_0_elements(157)); -- 
    -- CP-element group 158:  transition  input  output  bypass 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	155 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	159 
    -- CP-element group 158:  members (6) 
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_sample_completed_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_update_start_
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/$exit
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Sample/ra
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/$entry
      -- CP-element group 158: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/cr
      -- 
    ra_1861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_0, ack => testConfigure_CP_0_elements(158)); -- 
    cr_1865_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1865_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(158), ack => RPIPE_ConvTranspose_input_pipe_700_inst_req_1); -- 
    -- CP-element group 159:  transition  input  output  bypass 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	158 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	160 
    -- CP-element group 159:  members (6) 
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_update_completed_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/$exit
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_700_Update/ca
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/rr
      -- 
    ca_1866_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 159_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_700_inst_ack_1, ack => testConfigure_CP_0_elements(159)); -- 
    rr_1874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(159), ack => type_cast_704_inst_req_0); -- 
    -- CP-element group 160:  transition  input  bypass 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: 	159 
    -- CP-element group 160: successors 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_sample_completed_
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/$exit
      -- CP-element group 160: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Sample/ra
      -- 
    ra_1875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 160_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_0, ack => testConfigure_CP_0_elements(160)); -- 
    -- CP-element group 161:  transition  input  bypass 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	295 
    -- CP-element group 161: successors 
    -- CP-element group 161: 	162 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_update_completed_
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/$exit
      -- CP-element group 161: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/ca
      -- 
    ca_1880_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_704_inst_ack_1, ack => testConfigure_CP_0_elements(161)); -- 
    -- CP-element group 162:  join  transition  output  bypass 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	129 
    -- CP-element group 162: 	133 
    -- CP-element group 162: 	137 
    -- CP-element group 162: 	141 
    -- CP-element group 162: 	145 
    -- CP-element group 162: 	149 
    -- CP-element group 162: 	153 
    -- CP-element group 162: 	157 
    -- CP-element group 162: 	161 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (9) 
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_sample_start_
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/$exit
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/split_req
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/ptr_deref_712_Split/split_ack
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/$entry
      -- CP-element group 162: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/rr
      -- 
    rr_1918_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1918_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(162), ack => ptr_deref_712_store_0_req_0); -- 
    testConfigure_cp_element_group_162: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_162"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(129) & testConfigure_CP_0_elements(133) & testConfigure_CP_0_elements(137) & testConfigure_CP_0_elements(141) & testConfigure_CP_0_elements(145) & testConfigure_CP_0_elements(149) & testConfigure_CP_0_elements(153) & testConfigure_CP_0_elements(157) & testConfigure_CP_0_elements(161);
      gj_testConfigure_cp_element_group_162 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(162), clk => clk, reset => reset); --
    end block;
    -- CP-element group 163:  transition  input  bypass 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	162 
    -- CP-element group 163: successors 
    -- CP-element group 163:  members (5) 
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_sample_completed_
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/$exit
      -- CP-element group 163: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Sample/word_access_start/word_0/ra
      -- 
    ra_1919_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 163_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_712_store_0_ack_0, ack => testConfigure_CP_0_elements(163)); -- 
    -- CP-element group 164:  transition  input  bypass 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: 	295 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	165 
    -- CP-element group 164:  members (5) 
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_update_completed_
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/$exit
      -- CP-element group 164: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/ca
      -- 
    ca_1930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 164_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_712_store_0_ack_1, ack => testConfigure_CP_0_elements(164)); -- 
    -- CP-element group 165:  branch  join  transition  place  output  bypass 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	126 
    -- CP-element group 165: 	164 
    -- CP-element group 165: successors 
    -- CP-element group 165: 	166 
    -- CP-element group 165: 	167 
    -- CP-element group 165:  members (10) 
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725__exit__
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726__entry__
      -- CP-element group 165: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_dead_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/$exit
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_eval_test/branch_req
      -- CP-element group 165: 	 branch_block_stmt_32/R_exitcond10_727_place
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_if_link/$entry
      -- CP-element group 165: 	 branch_block_stmt_32/if_stmt_726_else_link/$entry
      -- 
    branch_req_1938_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1938_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(165), ack => if_stmt_726_branch_req_0); -- 
    testConfigure_cp_element_group_165: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_165"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(126) & testConfigure_CP_0_elements(164);
      gj_testConfigure_cp_element_group_165 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(165), clk => clk, reset => reset); --
    end block;
    -- CP-element group 166:  merge  transition  place  input  bypass 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	165 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	289 
    -- CP-element group 166:  members (13) 
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506__exit__
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_726_if_link/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/if_stmt_726_if_link/if_choice_transition
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xbody67_forx_xcond119x_xpreheaderx_xloopexit_PhiReq/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiReqMerge
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/$exit
      -- CP-element group 166: 	 branch_block_stmt_32/merge_stmt_506_PhiAck/dummy
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$entry
      -- CP-element group 166: 	 branch_block_stmt_32/forx_xcond119x_xpreheaderx_xloopexit_forx_xcond119x_xpreheader_PhiReq/$exit
      -- 
    if_choice_transition_1943_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_726_branch_ack_1, ack => testConfigure_CP_0_elements(166)); -- 
    -- CP-element group 167:  fork  transition  place  input  output  bypass 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	165 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	291 
    -- CP-element group 167: 	292 
    -- CP-element group 167:  members (12) 
      -- CP-element group 167: 	 branch_block_stmt_32/if_stmt_726_else_link/$exit
      -- CP-element group 167: 	 branch_block_stmt_32/if_stmt_726_else_link/else_choice_transition
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/rr
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/$entry
      -- CP-element group 167: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/cr
      -- 
    else_choice_transition_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 167_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_726_branch_ack_0, ack => testConfigure_CP_0_elements(167)); -- 
    rr_3091_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3091_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_569_inst_req_0); -- 
    cr_3096_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3096_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(167), ack => type_cast_569_inst_req_1); -- 
    -- CP-element group 168:  transition  input  bypass 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: 	123 
    -- CP-element group 168: successors 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_sample_completed_
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/$exit
      -- CP-element group 168: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Sample/ra
      -- 
    ra_1961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 168_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_0, ack => testConfigure_CP_0_elements(168)); -- 
    -- CP-element group 169:  transition  place  input  bypass 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	123 
    -- CP-element group 169: successors 
    -- CP-element group 169: 	296 
    -- CP-element group 169:  members (9) 
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770__exit__
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_update_completed_
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/$exit
      -- CP-element group 169: 	 branch_block_stmt_32/assign_stmt_737_to_assign_stmt_770/type_cast_750_Update/ca
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/$entry
      -- CP-element group 169: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$entry
      -- 
    ca_1966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_750_inst_ack_1, ack => testConfigure_CP_0_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	301 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	209 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_sample_complete
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/$exit
      -- CP-element group 170: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/ack
      -- 
    ack_1995_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_785_index_offset_ack_0, ack => testConfigure_CP_0_elements(170)); -- 
    -- CP-element group 171:  transition  input  output  bypass 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	301 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (11) 
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_root_address_calculated
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_offset_calculated
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/$entry
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/$exit
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/sum_rename_req
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_base_plus_offset/sum_rename_ack
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/$entry
      -- CP-element group 171: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/req
      -- 
    ack_2000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 171_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_785_index_offset_ack_1, ack => testConfigure_CP_0_elements(171)); -- 
    req_2009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(171), ack => addr_of_786_final_reg_req_0); -- 
    -- CP-element group 172:  transition  input  bypass 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/$exit
      -- CP-element group 172: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_request/ack
      -- 
    ack_2010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_786_final_reg_ack_0, ack => testConfigure_CP_0_elements(172)); -- 
    -- CP-element group 173:  fork  transition  input  bypass 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	301 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	206 
    -- CP-element group 173:  members (19) 
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/root_register_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/root_register_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_addrgen/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/sum_rename_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/sum_rename_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_plus_offset/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/base_resize_ack
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/base_resize_req
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_addr_resize/$entry
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_address_resized
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_root_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_word_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_base_address_calculated
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/$exit
      -- CP-element group 173: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/ack
      -- 
    ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_786_final_reg_ack_1, ack => testConfigure_CP_0_elements(173)); -- 
    -- CP-element group 174:  transition  input  output  bypass 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	301 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	175 
    -- CP-element group 174:  members (6) 
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_sample_completed_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_update_start_
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/$exit
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/ra
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/$entry
      -- CP-element group 174: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/cr
      -- 
    ra_2024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_0, ack => testConfigure_CP_0_elements(174)); -- 
    cr_2028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(174), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_1); -- 
    -- CP-element group 175:  fork  transition  input  output  bypass 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	174 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	176 
    -- CP-element group 175: 	178 
    -- CP-element group 175:  members (9) 
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_update_completed_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/$exit
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Update/ca
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/rr
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_sample_start_
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/rr
      -- 
    ca_2029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 175_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_789_inst_ack_1, ack => testConfigure_CP_0_elements(175)); -- 
    rr_2037_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2037_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => type_cast_793_inst_req_0); -- 
    rr_2051_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2051_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(175), ack => RPIPE_ConvTranspose_input_pipe_802_inst_req_0); -- 
    -- CP-element group 176:  transition  input  bypass 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	175 
    -- CP-element group 176: successors 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_sample_completed_
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/$exit
      -- CP-element group 176: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Sample/ra
      -- 
    ra_2038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 176_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_0, ack => testConfigure_CP_0_elements(176)); -- 
    -- CP-element group 177:  transition  input  bypass 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	301 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	206 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_update_completed_
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/$exit
      -- CP-element group 177: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/ca
      -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_793_inst_ack_1, ack => testConfigure_CP_0_elements(177)); -- 
    -- CP-element group 178:  transition  input  output  bypass 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	175 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	179 
    -- CP-element group 178:  members (6) 
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_sample_completed_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_update_start_
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/$exit
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Sample/ra
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/$entry
      -- CP-element group 178: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/cr
      -- 
    ra_2052_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_802_inst_ack_0, ack => testConfigure_CP_0_elements(178)); -- 
    cr_2056_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2056_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(178), ack => RPIPE_ConvTranspose_input_pipe_802_inst_req_1); -- 
    -- CP-element group 179:  fork  transition  input  output  bypass 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	178 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	180 
    -- CP-element group 179: 	182 
    -- CP-element group 179:  members (9) 
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_update_completed_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/$exit
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_802_Update/ca
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/rr
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_sample_start_
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/rr
      -- 
    ca_2057_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 179_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_802_inst_ack_1, ack => testConfigure_CP_0_elements(179)); -- 
    rr_2065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => type_cast_806_inst_req_0); -- 
    rr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(179), ack => RPIPE_ConvTranspose_input_pipe_820_inst_req_0); -- 
    -- CP-element group 180:  transition  input  bypass 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	179 
    -- CP-element group 180: successors 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_sample_completed_
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/$exit
      -- CP-element group 180: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Sample/ra
      -- 
    ra_2066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 180_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_0, ack => testConfigure_CP_0_elements(180)); -- 
    -- CP-element group 181:  transition  input  bypass 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	301 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	206 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_update_completed_
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/$exit
      -- CP-element group 181: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/ca
      -- 
    ca_2071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_806_inst_ack_1, ack => testConfigure_CP_0_elements(181)); -- 
    -- CP-element group 182:  transition  input  output  bypass 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	179 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (6) 
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_sample_completed_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_update_start_
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/$exit
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Sample/ra
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/$entry
      -- CP-element group 182: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/cr
      -- 
    ra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_820_inst_ack_0, ack => testConfigure_CP_0_elements(182)); -- 
    cr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(182), ack => RPIPE_ConvTranspose_input_pipe_820_inst_req_1); -- 
    -- CP-element group 183:  fork  transition  input  output  bypass 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	182 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	184 
    -- CP-element group 183: 	186 
    -- CP-element group 183:  members (9) 
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_update_completed_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/$exit
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_820_Update/ca
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/rr
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/$entry
      -- CP-element group 183: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/rr
      -- 
    ca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_820_inst_ack_1, ack => testConfigure_CP_0_elements(183)); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => type_cast_824_inst_req_0); -- 
    rr_2107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(183), ack => RPIPE_ConvTranspose_input_pipe_838_inst_req_0); -- 
    -- CP-element group 184:  transition  input  bypass 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	183 
    -- CP-element group 184: successors 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_sample_completed_
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/$exit
      -- CP-element group 184: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Sample/ra
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 184_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_0, ack => testConfigure_CP_0_elements(184)); -- 
    -- CP-element group 185:  transition  input  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	301 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	206 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_update_completed_
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/ca
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_824_inst_ack_1, ack => testConfigure_CP_0_elements(185)); -- 
    -- CP-element group 186:  transition  input  output  bypass 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	183 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	187 
    -- CP-element group 186:  members (6) 
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_sample_completed_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_update_start_
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/$exit
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Sample/ra
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/$entry
      -- CP-element group 186: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/cr
      -- 
    ra_2108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_838_inst_ack_0, ack => testConfigure_CP_0_elements(186)); -- 
    cr_2112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(186), ack => RPIPE_ConvTranspose_input_pipe_838_inst_req_1); -- 
    -- CP-element group 187:  fork  transition  input  output  bypass 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	186 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	188 
    -- CP-element group 187: 	190 
    -- CP-element group 187:  members (9) 
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/rr
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_update_completed_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/$exit
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_838_Update/ca
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_sample_start_
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/rr
      -- 
    ca_2113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 187_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_838_inst_ack_1, ack => testConfigure_CP_0_elements(187)); -- 
    rr_2121_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2121_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => type_cast_842_inst_req_0); -- 
    rr_2135_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2135_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(187), ack => RPIPE_ConvTranspose_input_pipe_856_inst_req_0); -- 
    -- CP-element group 188:  transition  input  bypass 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: 	187 
    -- CP-element group 188: successors 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_sample_completed_
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/$exit
      -- CP-element group 188: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Sample/ra
      -- 
    ra_2122_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 188_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_0, ack => testConfigure_CP_0_elements(188)); -- 
    -- CP-element group 189:  transition  input  bypass 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	301 
    -- CP-element group 189: successors 
    -- CP-element group 189: 	206 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/ca
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/$exit
      -- CP-element group 189: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_update_completed_
      -- 
    ca_2127_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_842_inst_ack_1, ack => testConfigure_CP_0_elements(189)); -- 
    -- CP-element group 190:  transition  input  output  bypass 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	187 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	191 
    -- CP-element group 190:  members (6) 
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_sample_completed_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/$exit
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/$entry
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_update_start_
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/cr
      -- CP-element group 190: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Sample/ra
      -- 
    ra_2136_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_856_inst_ack_0, ack => testConfigure_CP_0_elements(190)); -- 
    cr_2140_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2140_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(190), ack => RPIPE_ConvTranspose_input_pipe_856_inst_req_1); -- 
    -- CP-element group 191:  fork  transition  input  output  bypass 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	190 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	192 
    -- CP-element group 191: 	194 
    -- CP-element group 191:  members (9) 
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/$exit
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_sample_start_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_update_completed_
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_856_Update/ca
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/rr
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_sample_start_
      -- 
    ca_2141_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 191_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_856_inst_ack_1, ack => testConfigure_CP_0_elements(191)); -- 
    rr_2149_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2149_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => type_cast_860_inst_req_0); -- 
    rr_2163_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2163_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(191), ack => RPIPE_ConvTranspose_input_pipe_874_inst_req_0); -- 
    -- CP-element group 192:  transition  input  bypass 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: 	191 
    -- CP-element group 192: successors 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_sample_completed_
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/$exit
      -- CP-element group 192: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Sample/ra
      -- 
    ra_2150_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 192_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_0, ack => testConfigure_CP_0_elements(192)); -- 
    -- CP-element group 193:  transition  input  bypass 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	301 
    -- CP-element group 193: successors 
    -- CP-element group 193: 	206 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_update_completed_
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/ca
      -- CP-element group 193: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/$exit
      -- 
    ca_2155_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_860_inst_ack_1, ack => testConfigure_CP_0_elements(193)); -- 
    -- CP-element group 194:  transition  input  output  bypass 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	191 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (6) 
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/cr
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/$entry
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/ra
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Sample/$exit
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_update_start_
      -- CP-element group 194: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_sample_completed_
      -- 
    ra_2164_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_874_inst_ack_0, ack => testConfigure_CP_0_elements(194)); -- 
    cr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2168_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(194), ack => RPIPE_ConvTranspose_input_pipe_874_inst_req_1); -- 
    -- CP-element group 195:  fork  transition  input  output  bypass 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195: 	198 
    -- CP-element group 195:  members (9) 
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_sample_start_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/$exit
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_Update/ca
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_874_update_completed_
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/rr
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_sample_start_
      -- 
    ca_2169_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 195_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_874_inst_ack_1, ack => testConfigure_CP_0_elements(195)); -- 
    rr_2177_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2177_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => type_cast_878_inst_req_0); -- 
    rr_2191_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2191_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(195), ack => RPIPE_ConvTranspose_input_pipe_892_inst_req_0); -- 
    -- CP-element group 196:  transition  input  bypass 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196:  members (3) 
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_sample_completed_
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Sample/ra
      -- 
    ra_2178_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_0, ack => testConfigure_CP_0_elements(196)); -- 
    -- CP-element group 197:  transition  input  bypass 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	301 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	206 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_update_completed_
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/ca
      -- 
    ca_2183_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_878_inst_ack_1, ack => testConfigure_CP_0_elements(197)); -- 
    -- CP-element group 198:  transition  input  output  bypass 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	195 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	199 
    -- CP-element group 198:  members (6) 
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/cr
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/$entry
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/ra
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Sample/$exit
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_update_start_
      -- CP-element group 198: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_sample_completed_
      -- 
    ra_2192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 198_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_892_inst_ack_0, ack => testConfigure_CP_0_elements(198)); -- 
    cr_2196_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2196_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(198), ack => RPIPE_ConvTranspose_input_pipe_892_inst_req_1); -- 
    -- CP-element group 199:  fork  transition  input  output  bypass 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: 	198 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	200 
    -- CP-element group 199: 	202 
    -- CP-element group 199:  members (9) 
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/rr
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/$entry
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_sample_start_
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/ca
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_Update/$exit
      -- CP-element group 199: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_892_update_completed_
      -- 
    ca_2197_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 199_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_892_inst_ack_1, ack => testConfigure_CP_0_elements(199)); -- 
    rr_2205_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2205_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => type_cast_896_inst_req_0); -- 
    rr_2219_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2219_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(199), ack => RPIPE_ConvTranspose_input_pipe_910_inst_req_0); -- 
    -- CP-element group 200:  transition  input  bypass 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	199 
    -- CP-element group 200: successors 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/ra
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Sample/$exit
      -- CP-element group 200: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_sample_completed_
      -- 
    ra_2206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_0, ack => testConfigure_CP_0_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	301 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	206 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/ca
      -- CP-element group 201: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_update_completed_
      -- 
    ca_2211_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_896_inst_ack_1, ack => testConfigure_CP_0_elements(201)); -- 
    -- CP-element group 202:  transition  input  output  bypass 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	199 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	203 
    -- CP-element group 202:  members (6) 
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_sample_completed_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_update_start_
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/$exit
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Sample/ra
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/$entry
      -- CP-element group 202: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/cr
      -- 
    ra_2220_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 202_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_910_inst_ack_0, ack => testConfigure_CP_0_elements(202)); -- 
    cr_2224_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2224_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(202), ack => RPIPE_ConvTranspose_input_pipe_910_inst_req_1); -- 
    -- CP-element group 203:  transition  input  output  bypass 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: 	202 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	204 
    -- CP-element group 203:  members (6) 
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/$entry
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_update_completed_
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/rr
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/$exit
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_910_Update/ca
      -- CP-element group 203: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_sample_start_
      -- 
    ca_2225_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 203_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_ConvTranspose_input_pipe_910_inst_ack_1, ack => testConfigure_CP_0_elements(203)); -- 
    rr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(203), ack => type_cast_914_inst_req_0); -- 
    -- CP-element group 204:  transition  input  bypass 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	203 
    -- CP-element group 204: successors 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Sample/ra
      -- CP-element group 204: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_sample_completed_
      -- 
    ra_2234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_0, ack => testConfigure_CP_0_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	301 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	206 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/ca
      -- CP-element group 205: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_update_completed_
      -- 
    ca_2239_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_914_inst_ack_1, ack => testConfigure_CP_0_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	173 
    -- CP-element group 206: 	177 
    -- CP-element group 206: 	181 
    -- CP-element group 206: 	185 
    -- CP-element group 206: 	189 
    -- CP-element group 206: 	193 
    -- CP-element group 206: 	197 
    -- CP-element group 206: 	201 
    -- CP-element group 206: 	205 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	207 
    -- CP-element group 206:  members (9) 
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/rr
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/split_ack
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/split_req
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/$exit
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/ptr_deref_922_Split/$entry
      -- CP-element group 206: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/$entry
      -- 
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(206), ack => ptr_deref_922_store_0_req_0); -- 
    testConfigure_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(173) & testConfigure_CP_0_elements(177) & testConfigure_CP_0_elements(181) & testConfigure_CP_0_elements(185) & testConfigure_CP_0_elements(189) & testConfigure_CP_0_elements(193) & testConfigure_CP_0_elements(197) & testConfigure_CP_0_elements(201) & testConfigure_CP_0_elements(205);
      gj_testConfigure_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  transition  input  bypass 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: 	206 
    -- CP-element group 207: successors 
    -- CP-element group 207:  members (5) 
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_sample_completed_
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/ra
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/word_0/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/word_access_start/$exit
      -- CP-element group 207: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Sample/$exit
      -- 
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 207_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_922_store_0_ack_0, ack => testConfigure_CP_0_elements(207)); -- 
    -- CP-element group 208:  transition  input  bypass 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	301 
    -- CP-element group 208: successors 
    -- CP-element group 208: 	209 
    -- CP-element group 208:  members (5) 
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/ca
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/$exit
      -- CP-element group 208: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_update_completed_
      -- 
    ca_2289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_922_store_0_ack_1, ack => testConfigure_CP_0_elements(208)); -- 
    -- CP-element group 209:  branch  join  transition  place  output  bypass 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	170 
    -- CP-element group 209: 	208 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	210 
    -- CP-element group 209: 	211 
    -- CP-element group 209:  members (10) 
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935__exit__
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936__entry__
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_else_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_if_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/branch_req
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/$exit
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_eval_test/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/if_stmt_936_dead_link/$entry
      -- CP-element group 209: 	 branch_block_stmt_32/R_exitcond19_937_place
      -- CP-element group 209: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/$exit
      -- 
    branch_req_2297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(209), ack => if_stmt_936_branch_req_0); -- 
    testConfigure_cp_element_group_209: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_209"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(170) & testConfigure_CP_0_elements(208);
      gj_testConfigure_cp_element_group_209 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(209), clk => clk, reset => reset); --
    end block;
    -- CP-element group 210:  merge  transition  place  input  bypass 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	209 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	302 
    -- CP-element group 210:  members (13) 
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942__exit__
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_936_if_link/if_choice_transition
      -- CP-element group 210: 	 branch_block_stmt_32/if_stmt_936_if_link/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xbody126_forx_xend180x_xloopexit_PhiReq/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiReqMerge
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/$exit
      -- CP-element group 210: 	 branch_block_stmt_32/merge_stmt_942_PhiAck/dummy
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180_PhiReq/$entry
      -- CP-element group 210: 	 branch_block_stmt_32/forx_xend180x_xloopexit_forx_xend180_PhiReq/$exit
      -- 
    if_choice_transition_2302_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 210_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_936_branch_ack_1, ack => testConfigure_CP_0_elements(210)); -- 
    -- CP-element group 211:  fork  transition  place  input  output  bypass 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: 	209 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	297 
    -- CP-element group 211: 	298 
    -- CP-element group 211:  members (12) 
      -- CP-element group 211: 	 branch_block_stmt_32/if_stmt_936_else_link/else_choice_transition
      -- CP-element group 211: 	 branch_block_stmt_32/if_stmt_936_else_link/$exit
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/rr
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 211_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_936_branch_ack_0, ack => testConfigure_CP_0_elements(211)); -- 
    rr_3145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_779_inst_req_0); -- 
    cr_3150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(211), ack => type_cast_779_inst_req_1); -- 
    -- CP-element group 212:  transition  input  bypass 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	303 
    -- CP-element group 212: successors 
    -- CP-element group 212:  members (5) 
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/word_0/$exit
      -- CP-element group 212: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/word_0/ra
      -- 
    ra_2345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_955_load_0_ack_0, ack => testConfigure_CP_0_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	303 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (9) 
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/ptr_deref_955_Merge/merge_ack
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/ptr_deref_955_Merge/merge_req
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/ptr_deref_955_Merge/$exit
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/ptr_deref_955_Merge/$entry
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/word_0/ca
      -- CP-element group 213: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/word_0/$exit
      -- 
    ca_2356_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_955_load_0_ack_1, ack => testConfigure_CP_0_elements(213)); -- 
    -- CP-element group 214:  transition  input  bypass 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	303 
    -- CP-element group 214: successors 
    -- CP-element group 214:  members (5) 
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_sample_completed_
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/word_0/ra
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/word_0/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/$exit
      -- CP-element group 214: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/$exit
      -- 
    ra_2395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 214_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_967_load_0_ack_0, ack => testConfigure_CP_0_elements(214)); -- 
    -- CP-element group 215:  transition  input  bypass 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: 	303 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	218 
    -- CP-element group 215:  members (9) 
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_update_completed_
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/ptr_deref_967_Merge/merge_ack
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/ptr_deref_967_Merge/merge_req
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/ptr_deref_967_Merge/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/ptr_deref_967_Merge/$entry
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/word_0/ca
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/word_0/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/$exit
      -- CP-element group 215: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/$exit
      -- 
    ca_2406_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 215_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_967_load_0_ack_1, ack => testConfigure_CP_0_elements(215)); -- 
    -- CP-element group 216:  transition  input  bypass 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	303 
    -- CP-element group 216: successors 
    -- CP-element group 216:  members (5) 
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/word_0/ra
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/word_0/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_sample_completed_
      -- 
    ra_2445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_979_load_0_ack_0, ack => testConfigure_CP_0_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	303 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (9) 
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/word_0/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/word_0/ca
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/ptr_deref_979_Merge/$entry
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/ptr_deref_979_Merge/$exit
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/ptr_deref_979_Merge/merge_req
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/ptr_deref_979_Merge/merge_ack
      -- CP-element group 217: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_update_completed_
      -- 
    ca_2456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_979_load_0_ack_1, ack => testConfigure_CP_0_elements(217)); -- 
    -- CP-element group 218:  branch  join  transition  place  output  bypass 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	215 
    -- CP-element group 218: 	217 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	219 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (10) 
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_else_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996__exit__
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997__entry__
      -- CP-element group 218: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_if_link/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/R_cmp191204_998_place
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_eval_test/branch_req
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_eval_test/$exit
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_eval_test/$entry
      -- CP-element group 218: 	 branch_block_stmt_32/if_stmt_997_dead_link/$entry
      -- 
    branch_req_2469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(218), ack => if_stmt_997_branch_req_0); -- 
    testConfigure_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(213) & testConfigure_CP_0_elements(215) & testConfigure_CP_0_elements(217);
      gj_testConfigure_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: 	218 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: 	222 
    -- CP-element group 219:  members (18) 
      -- CP-element group 219: 	 branch_block_stmt_32/merge_stmt_1003__exit__
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038__entry__
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend180_bbx_xnph
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_sample_start_
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_997_if_link/if_choice_transition
      -- CP-element group 219: 	 branch_block_stmt_32/if_stmt_997_if_link/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Update/cr
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Sample/rr
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Sample/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_update_start_
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend180_bbx_xnph_PhiReq/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/forx_xend180_bbx_xnph_PhiReq/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/merge_stmt_1003_PhiReqMerge
      -- CP-element group 219: 	 branch_block_stmt_32/merge_stmt_1003_PhiAck/$entry
      -- CP-element group 219: 	 branch_block_stmt_32/merge_stmt_1003_PhiAck/$exit
      -- CP-element group 219: 	 branch_block_stmt_32/merge_stmt_1003_PhiAck/dummy
      -- 
    if_choice_transition_2474_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 219_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_997_branch_ack_1, ack => testConfigure_CP_0_elements(219)); -- 
    cr_2496_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2496_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1024_inst_req_1); -- 
    rr_2491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(219), ack => type_cast_1024_inst_req_0); -- 
    -- CP-element group 220:  transition  place  input  bypass 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: 	310 
    -- CP-element group 220:  members (5) 
      -- CP-element group 220: 	 branch_block_stmt_32/forx_xend180_forx_xend200
      -- CP-element group 220: 	 branch_block_stmt_32/if_stmt_997_else_link/else_choice_transition
      -- CP-element group 220: 	 branch_block_stmt_32/if_stmt_997_else_link/$exit
      -- CP-element group 220: 	 branch_block_stmt_32/forx_xend180_forx_xend200_PhiReq/$entry
      -- CP-element group 220: 	 branch_block_stmt_32/forx_xend180_forx_xend200_PhiReq/$exit
      -- 
    else_choice_transition_2478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_997_branch_ack_0, ack => testConfigure_CP_0_elements(220)); -- 
    -- CP-element group 221:  transition  input  bypass 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_sample_completed_
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Sample/ra
      -- CP-element group 221: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Sample/$exit
      -- 
    ra_2492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1024_inst_ack_0, ack => testConfigure_CP_0_elements(221)); -- 
    -- CP-element group 222:  transition  place  input  bypass 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	219 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	304 
    -- CP-element group 222:  members (9) 
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038__exit__
      -- CP-element group 222: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Update/ca
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_Update/$exit
      -- CP-element group 222: 	 branch_block_stmt_32/assign_stmt_1009_to_assign_stmt_1038/type_cast_1024_update_completed_
      -- CP-element group 222: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/$entry
      -- CP-element group 222: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$entry
      -- 
    ca_2497_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 222_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1024_inst_ack_1, ack => testConfigure_CP_0_elements(222)); -- 
    -- CP-element group 223:  transition  input  bypass 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	309 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	229 
    -- CP-element group 223:  members (3) 
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Sample/ack
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Sample/$exit
      -- CP-element group 223: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_sample_complete
      -- 
    ack_2526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 223_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_index_offset_ack_0, ack => testConfigure_CP_0_elements(223)); -- 
    -- CP-element group 224:  transition  input  output  bypass 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	309 
    -- CP-element group 224: successors 
    -- CP-element group 224: 	225 
    -- CP-element group 224:  members (11) 
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Update/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_root_address_calculated
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Update/ack
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_offset_calculated
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_request/req
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_request/$entry
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_base_plus_offset/sum_rename_ack
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_base_plus_offset/sum_rename_req
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_base_plus_offset/$exit
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_base_plus_offset/$entry
      -- CP-element group 224: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_sample_start_
      -- 
    ack_2531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1053_index_offset_ack_1, ack => testConfigure_CP_0_elements(224)); -- 
    req_2540_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2540_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(224), ack => addr_of_1054_final_reg_req_0); -- 
    -- CP-element group 225:  transition  input  bypass 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	224 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (3) 
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_request/ack
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_sample_completed_
      -- CP-element group 225: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_request/$exit
      -- 
    ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1054_final_reg_ack_0, ack => testConfigure_CP_0_elements(225)); -- 
    -- CP-element group 226:  join  fork  transition  input  output  bypass 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	309 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	227 
    -- CP-element group 226:  members (28) 
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_complete/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_plus_offset/sum_rename_ack
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_complete/ack
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_update_completed_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_addr_resize/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_plus_offset/sum_rename_req
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_address_resized
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_plus_offset/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_root_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_word_address_calculated
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_word_addrgen/root_register_ack
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_sample_start_
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_plus_offset/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_word_addrgen/root_register_req
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_word_addrgen/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/word_0/rr
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/ptr_deref_1057_Split/split_ack
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_word_addrgen/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/word_0/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/ptr_deref_1057_Split/split_req
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/ptr_deref_1057_Split/$entry
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/ptr_deref_1057_Split/$exit
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_addr_resize/base_resize_ack
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_addr_resize/base_resize_req
      -- CP-element group 226: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_base_addr_resize/$exit
      -- 
    ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 226_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1054_final_reg_ack_1, ack => testConfigure_CP_0_elements(226)); -- 
    rr_2584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(226), ack => ptr_deref_1057_store_0_req_0); -- 
    -- CP-element group 227:  transition  input  bypass 
    -- CP-element group 227: predecessors 
    -- CP-element group 227: 	226 
    -- CP-element group 227: successors 
    -- CP-element group 227:  members (5) 
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_sample_completed_
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/$exit
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/word_0/ra
      -- CP-element group 227: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Sample/word_access_start/word_0/$exit
      -- 
    ra_2585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 227_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1057_store_0_ack_0, ack => testConfigure_CP_0_elements(227)); -- 
    -- CP-element group 228:  transition  input  bypass 
    -- CP-element group 228: predecessors 
    -- CP-element group 228: 	309 
    -- CP-element group 228: successors 
    -- CP-element group 228: 	229 
    -- CP-element group 228:  members (5) 
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_update_completed_
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/word_0/$exit
      -- CP-element group 228: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/word_0/ca
      -- 
    ca_2596_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 228_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1057_store_0_ack_1, ack => testConfigure_CP_0_elements(228)); -- 
    -- CP-element group 229:  branch  join  transition  place  output  bypass 
    -- CP-element group 229: predecessors 
    -- CP-element group 229: 	223 
    -- CP-element group 229: 	228 
    -- CP-element group 229: successors 
    -- CP-element group 229: 	230 
    -- CP-element group 229: 	231 
    -- CP-element group 229:  members (10) 
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071__exit__
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072__entry__
      -- CP-element group 229: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_dead_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_eval_test/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_eval_test/$exit
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_eval_test/branch_req
      -- CP-element group 229: 	 branch_block_stmt_32/R_exitcond20_1073_place
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_if_link/$entry
      -- CP-element group 229: 	 branch_block_stmt_32/if_stmt_1072_else_link/$entry
      -- 
    branch_req_2604_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2604_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(229), ack => if_stmt_1072_branch_req_0); -- 
    testConfigure_cp_element_group_229: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_229"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(223) & testConfigure_CP_0_elements(228);
      gj_testConfigure_cp_element_group_229 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(229), clk => clk, reset => reset); --
    end block;
    -- CP-element group 230:  merge  transition  place  input  bypass 
    -- CP-element group 230: predecessors 
    -- CP-element group 230: 	229 
    -- CP-element group 230: successors 
    -- CP-element group 230: 	310 
    -- CP-element group 230:  members (13) 
      -- CP-element group 230: 	 branch_block_stmt_32/merge_stmt_1078__exit__
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xend200x_xloopexit_forx_xend200
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_1072_if_link/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/if_stmt_1072_if_link/if_choice_transition
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody193_forx_xend200x_xloopexit
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xbody193_forx_xend200x_xloopexit_PhiReq/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/merge_stmt_1078_PhiReqMerge
      -- CP-element group 230: 	 branch_block_stmt_32/merge_stmt_1078_PhiAck/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/merge_stmt_1078_PhiAck/$exit
      -- CP-element group 230: 	 branch_block_stmt_32/merge_stmt_1078_PhiAck/dummy
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xend200x_xloopexit_forx_xend200_PhiReq/$entry
      -- CP-element group 230: 	 branch_block_stmt_32/forx_xend200x_xloopexit_forx_xend200_PhiReq/$exit
      -- 
    if_choice_transition_2609_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 230_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1072_branch_ack_1, ack => testConfigure_CP_0_elements(230)); -- 
    -- CP-element group 231:  fork  transition  place  input  output  bypass 
    -- CP-element group 231: predecessors 
    -- CP-element group 231: 	229 
    -- CP-element group 231: successors 
    -- CP-element group 231: 	305 
    -- CP-element group 231: 	306 
    -- CP-element group 231:  members (12) 
      -- CP-element group 231: 	 branch_block_stmt_32/if_stmt_1072_else_link/$exit
      -- CP-element group 231: 	 branch_block_stmt_32/if_stmt_1072_else_link/else_choice_transition
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Sample/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Sample/rr
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Update/$entry
      -- CP-element group 231: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Update/cr
      -- 
    else_choice_transition_2613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 231_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1072_branch_ack_0, ack => testConfigure_CP_0_elements(231)); -- 
    rr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1047_inst_req_0); -- 
    cr_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(231), ack => type_cast_1047_inst_req_1); -- 
    -- CP-element group 232:  transition  input  bypass 
    -- CP-element group 232: predecessors 
    -- CP-element group 232: 	310 
    -- CP-element group 232: successors 
    -- CP-element group 232:  members (3) 
      -- CP-element group 232: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_sample_completed_
      -- CP-element group 232: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Sample/$exit
      -- CP-element group 232: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Sample/ra
      -- 
    ra_2627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 232_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_0, ack => testConfigure_CP_0_elements(232)); -- 
    -- CP-element group 233:  transition  place  input  bypass 
    -- CP-element group 233: predecessors 
    -- CP-element group 233: 	310 
    -- CP-element group 233: successors 
    -- CP-element group 233:  members (16) 
      -- CP-element group 233: 	 $exit
      -- CP-element group 233: 	 branch_block_stmt_32/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/branch_block_stmt_32__exit__
      -- CP-element group 233: 	 branch_block_stmt_32/assign_stmt_1084__exit__
      -- CP-element group 233: 	 branch_block_stmt_32/return__
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_1086__exit__
      -- CP-element group 233: 	 branch_block_stmt_32/assign_stmt_1084/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_update_completed_
      -- CP-element group 233: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Update/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Update/ca
      -- CP-element group 233: 	 branch_block_stmt_32/return___PhiReq/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/return___PhiReq/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_1086_PhiReqMerge
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_1086_PhiAck/$entry
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_1086_PhiAck/$exit
      -- CP-element group 233: 	 branch_block_stmt_32/merge_stmt_1086_PhiAck/dummy
      -- 
    ca_2632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 233_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1083_inst_ack_1, ack => testConfigure_CP_0_elements(233)); -- 
    -- CP-element group 234:  transition  input  bypass 
    -- CP-element group 234: predecessors 
    -- CP-element group 234: 	32 
    -- CP-element group 234: successors 
    -- CP-element group 234: 	236 
    -- CP-element group 234:  members (2) 
      -- CP-element group 234: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/$exit
      -- CP-element group 234: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Sample/ra
      -- 
    ra_2664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 234_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_0, ack => testConfigure_CP_0_elements(234)); -- 
    -- CP-element group 235:  transition  input  bypass 
    -- CP-element group 235: predecessors 
    -- CP-element group 235: 	32 
    -- CP-element group 235: successors 
    -- CP-element group 235: 	236 
    -- CP-element group 235:  members (2) 
      -- CP-element group 235: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/$exit
      -- CP-element group 235: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/Update/ca
      -- 
    ca_2669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 235_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_76_inst_ack_1, ack => testConfigure_CP_0_elements(235)); -- 
    -- CP-element group 236:  join  transition  output  bypass 
    -- CP-element group 236: predecessors 
    -- CP-element group 236: 	234 
    -- CP-element group 236: 	235 
    -- CP-element group 236: successors 
    -- CP-element group 236: 	240 
    -- CP-element group 236:  members (5) 
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_76/SplitProtocol/$exit
      -- CP-element group 236: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- 
    phi_stmt_73_req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2670_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(236), ack => phi_stmt_73_req_0); -- 
    testConfigure_cp_element_group_236: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_236"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(234) & testConfigure_CP_0_elements(235);
      gj_testConfigure_cp_element_group_236 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(236), clk => clk, reset => reset); --
    end block;
    -- CP-element group 237:  transition  input  bypass 
    -- CP-element group 237: predecessors 
    -- CP-element group 237: 	32 
    -- CP-element group 237: successors 
    -- CP-element group 237: 	239 
    -- CP-element group 237:  members (2) 
      -- CP-element group 237: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/$exit
      -- CP-element group 237: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Sample/ra
      -- 
    ra_2687_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 237_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_0, ack => testConfigure_CP_0_elements(237)); -- 
    -- CP-element group 238:  transition  input  bypass 
    -- CP-element group 238: predecessors 
    -- CP-element group 238: 	32 
    -- CP-element group 238: successors 
    -- CP-element group 238: 	239 
    -- CP-element group 238:  members (2) 
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/$exit
      -- CP-element group 238: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/Update/ca
      -- 
    ca_2692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 238_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_83_inst_ack_1, ack => testConfigure_CP_0_elements(238)); -- 
    -- CP-element group 239:  join  transition  output  bypass 
    -- CP-element group 239: predecessors 
    -- CP-element group 239: 	237 
    -- CP-element group 239: 	238 
    -- CP-element group 239: successors 
    -- CP-element group 239: 	240 
    -- CP-element group 239:  members (5) 
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_83/SplitProtocol/$exit
      -- CP-element group 239: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2693_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2693_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(239), ack => phi_stmt_80_req_0); -- 
    testConfigure_cp_element_group_239: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_239"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(237) & testConfigure_CP_0_elements(238);
      gj_testConfigure_cp_element_group_239 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(239), clk => clk, reset => reset); --
    end block;
    -- CP-element group 240:  join  transition  bypass 
    -- CP-element group 240: predecessors 
    -- CP-element group 240: 	236 
    -- CP-element group 240: 	239 
    -- CP-element group 240: successors 
    -- CP-element group 240: 	246 
    -- CP-element group 240:  members (1) 
      -- CP-element group 240: 	 branch_block_stmt_32/forx_xbody_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_240: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_240"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(236) & testConfigure_CP_0_elements(239);
      gj_testConfigure_cp_element_group_240 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(240), clk => clk, reset => reset); --
    end block;
    -- CP-element group 241:  transition  output  delay-element  bypass 
    -- CP-element group 241: predecessors 
    -- CP-element group 241: 	14 
    -- CP-element group 241: successors 
    -- CP-element group 241: 	245 
    -- CP-element group 241:  members (4) 
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/$exit
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_sources/type_cast_79_konst_delay_trans
      -- CP-element group 241: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_73/phi_stmt_73_req
      -- 
    phi_stmt_73_req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_73_req_2704_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(241), ack => phi_stmt_73_req_1); -- 
    -- Element group testConfigure_CP_0_elements(241) is a control-delay.
    cp_element_241_delay: control_delay_element  generic map(name => " 241_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(14), ack => testConfigure_CP_0_elements(241), clk => clk, reset =>reset);
    -- CP-element group 242:  transition  input  bypass 
    -- CP-element group 242: predecessors 
    -- CP-element group 242: 	14 
    -- CP-element group 242: successors 
    -- CP-element group 242: 	244 
    -- CP-element group 242:  members (2) 
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/$exit
      -- CP-element group 242: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Sample/ra
      -- 
    ra_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 242_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_0, ack => testConfigure_CP_0_elements(242)); -- 
    -- CP-element group 243:  transition  input  bypass 
    -- CP-element group 243: predecessors 
    -- CP-element group 243: 	14 
    -- CP-element group 243: successors 
    -- CP-element group 243: 	244 
    -- CP-element group 243:  members (2) 
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/$exit
      -- CP-element group 243: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/Update/ca
      -- 
    ca_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 243_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_85_inst_ack_1, ack => testConfigure_CP_0_elements(243)); -- 
    -- CP-element group 244:  join  transition  output  bypass 
    -- CP-element group 244: predecessors 
    -- CP-element group 244: 	242 
    -- CP-element group 244: 	243 
    -- CP-element group 244: successors 
    -- CP-element group 244: 	245 
    -- CP-element group 244:  members (5) 
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_sources/type_cast_85/SplitProtocol/$exit
      -- CP-element group 244: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/phi_stmt_80/phi_stmt_80_req
      -- 
    phi_stmt_80_req_2727_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_80_req_2727_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(244), ack => phi_stmt_80_req_1); -- 
    testConfigure_cp_element_group_244: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_244"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(242) & testConfigure_CP_0_elements(243);
      gj_testConfigure_cp_element_group_244 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(244), clk => clk, reset => reset); --
    end block;
    -- CP-element group 245:  join  transition  bypass 
    -- CP-element group 245: predecessors 
    -- CP-element group 245: 	241 
    -- CP-element group 245: 	244 
    -- CP-element group 245: successors 
    -- CP-element group 245: 	246 
    -- CP-element group 245:  members (1) 
      -- CP-element group 245: 	 branch_block_stmt_32/forx_xbodyx_xpreheader_forx_xbody_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_245: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_245"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(241) & testConfigure_CP_0_elements(244);
      gj_testConfigure_cp_element_group_245 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(245), clk => clk, reset => reset); --
    end block;
    -- CP-element group 246:  merge  fork  transition  place  bypass 
    -- CP-element group 246: predecessors 
    -- CP-element group 246: 	240 
    -- CP-element group 246: 	245 
    -- CP-element group 246: successors 
    -- CP-element group 246: 	247 
    -- CP-element group 246: 	248 
    -- CP-element group 246:  members (2) 
      -- CP-element group 246: 	 branch_block_stmt_32/merge_stmt_72_PhiReqMerge
      -- CP-element group 246: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(246) <= OrReduce(testConfigure_CP_0_elements(240) & testConfigure_CP_0_elements(245));
    -- CP-element group 247:  transition  input  bypass 
    -- CP-element group 247: predecessors 
    -- CP-element group 247: 	246 
    -- CP-element group 247: successors 
    -- CP-element group 247: 	249 
    -- CP-element group 247:  members (1) 
      -- CP-element group 247: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_73_ack
      -- 
    phi_stmt_73_ack_2732_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 247_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_73_ack_0, ack => testConfigure_CP_0_elements(247)); -- 
    -- CP-element group 248:  transition  input  bypass 
    -- CP-element group 248: predecessors 
    -- CP-element group 248: 	246 
    -- CP-element group 248: successors 
    -- CP-element group 248: 	249 
    -- CP-element group 248:  members (1) 
      -- CP-element group 248: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/phi_stmt_80_ack
      -- 
    phi_stmt_80_ack_2733_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 248_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_80_ack_0, ack => testConfigure_CP_0_elements(248)); -- 
    -- CP-element group 249:  join  fork  transition  place  output  bypass 
    -- CP-element group 249: predecessors 
    -- CP-element group 249: 	247 
    -- CP-element group 249: 	248 
    -- CP-element group 249: successors 
    -- CP-element group 249: 	15 
    -- CP-element group 249: 	16 
    -- CP-element group 249: 	17 
    -- CP-element group 249: 	18 
    -- CP-element group 249: 	20 
    -- CP-element group 249: 	22 
    -- CP-element group 249: 	23 
    -- CP-element group 249: 	25 
    -- CP-element group 249: 	26 
    -- CP-element group 249: 	29 
    -- CP-element group 249:  members (61) 
      -- CP-element group 249: 	 branch_block_stmt_32/merge_stmt_72__exit__
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135__entry__
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_root_address_calculated
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_address_resized
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/base_resize_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_addr_resize/base_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_95_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resized_1
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scaled_1
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_computed_1
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/index_resize_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_resize_1/index_resize_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/scale_rename_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_index_scale_1/scale_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_update_start
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Sample/req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/array_obj_ref_101_final_index_sum_regn_Update/req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/addr_of_102_complete/req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_105_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/sum_rename_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_base_plus_offset/sum_rename_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/$exit
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/root_register_req
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_word_addrgen/root_register_ack
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/ptr_deref_122_Update/word_access_complete/word_0/cr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_sample_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/RPIPE_ConvTranspose_input_pipe_130_Sample/rr
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_update_start_
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/$entry
      -- CP-element group 249: 	 branch_block_stmt_32/assign_stmt_92_to_assign_stmt_135/type_cast_134_Update/cr
      -- CP-element group 249: 	 branch_block_stmt_32/merge_stmt_72_PhiAck/$exit
      -- 
    rr_246_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_246_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_95_inst_req_0); -- 
    cr_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_95_inst_req_1); -- 
    req_277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_101_index_offset_req_0); -- 
    req_282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => array_obj_ref_101_index_offset_req_1); -- 
    req_297_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_297_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => addr_of_102_final_reg_req_1); -- 
    cr_347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_105_store_0_req_1); -- 
    cr_392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => ptr_deref_122_load_0_req_1); -- 
    rr_406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => RPIPE_ConvTranspose_input_pipe_130_inst_req_0); -- 
    cr_425_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_425_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(249), ack => type_cast_134_inst_req_1); -- 
    testConfigure_cp_element_group_249: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_249"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(247) & testConfigure_CP_0_elements(248);
      gj_testConfigure_cp_element_group_249 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(249), clk => clk, reset => reset); --
    end block;
    -- CP-element group 250:  transition  input  bypass 
    -- CP-element group 250: predecessors 
    -- CP-element group 250: 	33 
    -- CP-element group 250: successors 
    -- CP-element group 250: 	252 
    -- CP-element group 250:  members (2) 
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/$exit
      -- CP-element group 250: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Sample/ra
      -- 
    ra_2757_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 250_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_0, ack => testConfigure_CP_0_elements(250)); -- 
    -- CP-element group 251:  transition  input  bypass 
    -- CP-element group 251: predecessors 
    -- CP-element group 251: 	33 
    -- CP-element group 251: successors 
    -- CP-element group 251: 	252 
    -- CP-element group 251:  members (2) 
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/$exit
      -- CP-element group 251: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/Update/ca
      -- 
    ca_2762_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 251_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_146_inst_ack_1, ack => testConfigure_CP_0_elements(251)); -- 
    -- CP-element group 252:  join  transition  place  output  bypass 
    -- CP-element group 252: predecessors 
    -- CP-element group 252: 	250 
    -- CP-element group 252: 	251 
    -- CP-element group 252: successors 
    -- CP-element group 252: 	253 
    -- CP-element group 252:  members (8) 
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_sources/type_cast_146/SplitProtocol/$exit
      -- CP-element group 252: 	 branch_block_stmt_32/forx_xbody_forx_xendx_xloopexit_PhiReq/phi_stmt_143/phi_stmt_143_req
      -- CP-element group 252: 	 branch_block_stmt_32/merge_stmt_142_PhiReqMerge
      -- CP-element group 252: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/$entry
      -- 
    phi_stmt_143_req_2763_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_143_req_2763_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(252), ack => phi_stmt_143_req_0); -- 
    testConfigure_cp_element_group_252: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_252"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(250) & testConfigure_CP_0_elements(251);
      gj_testConfigure_cp_element_group_252 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(252), clk => clk, reset => reset); --
    end block;
    -- CP-element group 253:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 253: predecessors 
    -- CP-element group 253: 	252 
    -- CP-element group 253: successors 
    -- CP-element group 253: 	257 
    -- CP-element group 253: 	258 
    -- CP-element group 253:  members (13) 
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_142__exit__
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/$exit
      -- CP-element group 253: 	 branch_block_stmt_32/merge_stmt_142_PhiAck/phi_stmt_143_ack
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/rr
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/$entry
      -- CP-element group 253: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/cr
      -- 
    phi_stmt_143_ack_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 253_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_143_ack_0, ack => testConfigure_CP_0_elements(253)); -- 
    rr_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_155_inst_req_0); -- 
    cr_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(253), ack => type_cast_155_inst_req_1); -- 
    -- CP-element group 254:  transition  input  bypass 
    -- CP-element group 254: predecessors 
    -- CP-element group 254: 	13 
    -- CP-element group 254: successors 
    -- CP-element group 254: 	256 
    -- CP-element group 254:  members (2) 
      -- CP-element group 254: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/$exit
      -- CP-element group 254: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Sample/ra
      -- 
    ra_2788_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 254_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_0, ack => testConfigure_CP_0_elements(254)); -- 
    -- CP-element group 255:  transition  input  bypass 
    -- CP-element group 255: predecessors 
    -- CP-element group 255: 	13 
    -- CP-element group 255: successors 
    -- CP-element group 255: 	256 
    -- CP-element group 255:  members (2) 
      -- CP-element group 255: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/$exit
      -- CP-element group 255: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/Update/ca
      -- 
    ca_2793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 255_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_153_inst_ack_1, ack => testConfigure_CP_0_elements(255)); -- 
    -- CP-element group 256:  join  transition  output  bypass 
    -- CP-element group 256: predecessors 
    -- CP-element group 256: 	254 
    -- CP-element group 256: 	255 
    -- CP-element group 256: successors 
    -- CP-element group 256: 	260 
    -- CP-element group 256:  members (6) 
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_153/SplitProtocol/$exit
      -- CP-element group 256: 	 branch_block_stmt_32/entry_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- 
    phi_stmt_150_req_2794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(256), ack => phi_stmt_150_req_0); -- 
    testConfigure_cp_element_group_256: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_256"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(254) & testConfigure_CP_0_elements(255);
      gj_testConfigure_cp_element_group_256 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(256), clk => clk, reset => reset); --
    end block;
    -- CP-element group 257:  transition  input  bypass 
    -- CP-element group 257: predecessors 
    -- CP-element group 257: 	253 
    -- CP-element group 257: successors 
    -- CP-element group 257: 	259 
    -- CP-element group 257:  members (2) 
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/$exit
      -- CP-element group 257: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Sample/ra
      -- 
    ra_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 257_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_0, ack => testConfigure_CP_0_elements(257)); -- 
    -- CP-element group 258:  transition  input  bypass 
    -- CP-element group 258: predecessors 
    -- CP-element group 258: 	253 
    -- CP-element group 258: successors 
    -- CP-element group 258: 	259 
    -- CP-element group 258:  members (2) 
      -- CP-element group 258: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/$exit
      -- CP-element group 258: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/Update/ca
      -- 
    ca_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 258_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_155_inst_ack_1, ack => testConfigure_CP_0_elements(258)); -- 
    -- CP-element group 259:  join  transition  output  bypass 
    -- CP-element group 259: predecessors 
    -- CP-element group 259: 	257 
    -- CP-element group 259: 	258 
    -- CP-element group 259: successors 
    -- CP-element group 259: 	260 
    -- CP-element group 259:  members (6) 
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_sources/type_cast_155/SplitProtocol/$exit
      -- CP-element group 259: 	 branch_block_stmt_32/forx_xendx_xloopexit_forx_xend_PhiReq/phi_stmt_150/phi_stmt_150_req
      -- 
    phi_stmt_150_req_2820_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_150_req_2820_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(259), ack => phi_stmt_150_req_1); -- 
    testConfigure_cp_element_group_259: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_259"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(257) & testConfigure_CP_0_elements(258);
      gj_testConfigure_cp_element_group_259 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(259), clk => clk, reset => reset); --
    end block;
    -- CP-element group 260:  merge  transition  place  bypass 
    -- CP-element group 260: predecessors 
    -- CP-element group 260: 	256 
    -- CP-element group 260: 	259 
    -- CP-element group 260: successors 
    -- CP-element group 260: 	261 
    -- CP-element group 260:  members (2) 
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_149_PhiReqMerge
      -- CP-element group 260: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(260) <= OrReduce(testConfigure_CP_0_elements(256) & testConfigure_CP_0_elements(259));
    -- CP-element group 261:  join  fork  transition  place  input  output  bypass 
    -- CP-element group 261: predecessors 
    -- CP-element group 261: 	260 
    -- CP-element group 261: successors 
    -- CP-element group 261: 	34 
    -- CP-element group 261: 	35 
    -- CP-element group 261:  members (35) 
      -- CP-element group 261: 	 branch_block_stmt_32/merge_stmt_149__exit__
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172__entry__
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_sample_start_
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_update_start_
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_root_address_calculated
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_address_resized
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/base_resize_req
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_addr_resize/base_resize_ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/sum_rename_req
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_base_plus_offset/sum_rename_ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/root_register_req
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_word_addrgen/root_register_ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/split_req
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/ptr_deref_164_Split/split_ack
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Sample/word_access_start/word_0/rr
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/$entry
      -- CP-element group 261: 	 branch_block_stmt_32/assign_stmt_162_to_assign_stmt_172/ptr_deref_164_Update/word_access_complete/word_0/cr
      -- CP-element group 261: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/$exit
      -- CP-element group 261: 	 branch_block_stmt_32/merge_stmt_149_PhiAck/phi_stmt_150_ack
      -- 
    phi_stmt_150_ack_2825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 261_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_150_ack_0, ack => testConfigure_CP_0_elements(261)); -- 
    rr_487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_164_store_0_req_0); -- 
    cr_498_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_498_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(261), ack => ptr_deref_164_store_0_req_1); -- 
    -- CP-element group 262:  transition  input  bypass 
    -- CP-element group 262: predecessors 
    -- CP-element group 262: 	56 
    -- CP-element group 262: successors 
    -- CP-element group 262: 	264 
    -- CP-element group 262:  members (2) 
      -- CP-element group 262: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/$exit
      -- CP-element group 262: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Sample/ra
      -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 262_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_0, ack => testConfigure_CP_0_elements(262)); -- 
    -- CP-element group 263:  transition  input  bypass 
    -- CP-element group 263: predecessors 
    -- CP-element group 263: 	56 
    -- CP-element group 263: successors 
    -- CP-element group 263: 	264 
    -- CP-element group 263:  members (2) 
      -- CP-element group 263: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/$exit
      -- CP-element group 263: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/Update/ca
      -- 
    ca_2862_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 263_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_185_inst_ack_1, ack => testConfigure_CP_0_elements(263)); -- 
    -- CP-element group 264:  join  transition  output  bypass 
    -- CP-element group 264: predecessors 
    -- CP-element group 264: 	262 
    -- CP-element group 264: 	263 
    -- CP-element group 264: successors 
    -- CP-element group 264: 	266 
    -- CP-element group 264:  members (6) 
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_185/SplitProtocol/$exit
      -- CP-element group 264: 	 branch_block_stmt_32/forx_xbody14_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_req
      -- 
    phi_stmt_182_req_2863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_182_req_2863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(264), ack => phi_stmt_182_req_0); -- 
    testConfigure_cp_element_group_264: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_264"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(262) & testConfigure_CP_0_elements(263);
      gj_testConfigure_cp_element_group_264 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(264), clk => clk, reset => reset); --
    end block;
    -- CP-element group 265:  transition  output  delay-element  bypass 
    -- CP-element group 265: predecessors 
    -- CP-element group 265: 	37 
    -- CP-element group 265: successors 
    -- CP-element group 265: 	266 
    -- CP-element group 265:  members (5) 
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/$exit
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_sources/type_cast_188_konst_delay_trans
      -- CP-element group 265: 	 branch_block_stmt_32/forx_xbody14x_xpreheader_forx_xbody14_PhiReq/phi_stmt_182/phi_stmt_182_req
      -- 
    phi_stmt_182_req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_182_req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(265), ack => phi_stmt_182_req_1); -- 
    -- Element group testConfigure_CP_0_elements(265) is a control-delay.
    cp_element_265_delay: control_delay_element  generic map(name => " 265_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(37), ack => testConfigure_CP_0_elements(265), clk => clk, reset =>reset);
    -- CP-element group 266:  merge  transition  place  bypass 
    -- CP-element group 266: predecessors 
    -- CP-element group 266: 	264 
    -- CP-element group 266: 	265 
    -- CP-element group 266: successors 
    -- CP-element group 266: 	267 
    -- CP-element group 266:  members (2) 
      -- CP-element group 266: 	 branch_block_stmt_32/merge_stmt_181_PhiReqMerge
      -- CP-element group 266: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(266) <= OrReduce(testConfigure_CP_0_elements(264) & testConfigure_CP_0_elements(265));
    -- CP-element group 267:  fork  transition  place  input  output  bypass 
    -- CP-element group 267: predecessors 
    -- CP-element group 267: 	266 
    -- CP-element group 267: successors 
    -- CP-element group 267: 	47 
    -- CP-element group 267: 	40 
    -- CP-element group 267: 	41 
    -- CP-element group 267: 	43 
    -- CP-element group 267: 	44 
    -- CP-element group 267: 	38 
    -- CP-element group 267: 	39 
    -- CP-element group 267: 	50 
    -- CP-element group 267: 	51 
    -- CP-element group 267: 	53 
    -- CP-element group 267:  members (62) 
      -- CP-element group 267: 	 branch_block_stmt_32/merge_stmt_181__exit__
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238__entry__
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_198_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resized_1
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scaled_1
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_computed_1
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/index_resize_req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_resize_1/index_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/scale_rename_req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_index_scale_1/scale_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_update_start
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Sample/req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/array_obj_ref_204_final_index_sum_regn_Update/req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/addr_of_205_complete/req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_sample_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/RPIPE_ConvTranspose_input_pipe_208_Sample/rr
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/type_cast_212_Update/cr
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_215_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_update_start_
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_root_address_calculated
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_address_resized
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/base_resize_req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_addr_resize/base_resize_ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/sum_rename_req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_base_plus_offset/sum_rename_ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/root_register_req
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_word_addrgen/root_register_ack
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/$entry
      -- CP-element group 267: 	 branch_block_stmt_32/assign_stmt_195_to_assign_stmt_238/ptr_deref_232_Update/word_access_complete/word_0/cr
      -- CP-element group 267: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/$exit
      -- CP-element group 267: 	 branch_block_stmt_32/merge_stmt_181_PhiAck/phi_stmt_182_ack
      -- 
    phi_stmt_182_ack_2879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 267_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_182_ack_0, ack => testConfigure_CP_0_elements(267)); -- 
    rr_529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_198_inst_req_0); -- 
    cr_534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_198_inst_req_1); -- 
    req_560_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_560_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_204_index_offset_req_0); -- 
    req_565_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_565_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => array_obj_ref_204_index_offset_req_1); -- 
    req_580_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_580_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => addr_of_205_final_reg_req_1); -- 
    rr_589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => RPIPE_ConvTranspose_input_pipe_208_inst_req_0); -- 
    cr_608_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_608_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => type_cast_212_inst_req_1); -- 
    cr_658_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_658_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_215_store_0_req_1); -- 
    cr_703_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_703_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(267), ack => ptr_deref_232_load_0_req_1); -- 
    -- CP-element group 268:  merge  fork  transition  place  output  bypass 
    -- CP-element group 268: predecessors 
    -- CP-element group 268: 	36 
    -- CP-element group 268: 	57 
    -- CP-element group 268: successors 
    -- CP-element group 268: 	58 
    -- CP-element group 268: 	61 
    -- CP-element group 268:  members (13) 
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_247__exit__
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254__entry__
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_sample_start_
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/RPIPE_ConvTranspose_input_pipe_249_Sample/rr
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_update_start_
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/assign_stmt_250_to_assign_stmt_254/type_cast_253_Update/cr
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_247_PhiReqMerge
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/$entry
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/$exit
      -- CP-element group 268: 	 branch_block_stmt_32/merge_stmt_247_PhiAck/dummy
      -- 
    rr_740_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_740_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => RPIPE_ConvTranspose_input_pipe_249_inst_req_0); -- 
    cr_759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(268), ack => type_cast_253_inst_req_1); -- 
    testConfigure_CP_0_elements(268) <= OrReduce(testConfigure_CP_0_elements(36) & testConfigure_CP_0_elements(57));
    -- CP-element group 269:  transition  output  delay-element  bypass 
    -- CP-element group 269: predecessors 
    -- CP-element group 269: 	61 
    -- CP-element group 269: successors 
    -- CP-element group 269: 	273 
    -- CP-element group 269:  members (4) 
      -- CP-element group 269: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 269: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_261_konst_delay_trans
      -- CP-element group 269: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- 
    phi_stmt_257_req_2913_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_2913_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(269), ack => phi_stmt_257_req_0); -- 
    -- Element group testConfigure_CP_0_elements(269) is a control-delay.
    cp_element_269_delay: control_delay_element  generic map(name => " 269_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(61), ack => testConfigure_CP_0_elements(269), clk => clk, reset =>reset);
    -- CP-element group 270:  transition  input  bypass 
    -- CP-element group 270: predecessors 
    -- CP-element group 270: 	61 
    -- CP-element group 270: successors 
    -- CP-element group 270: 	272 
    -- CP-element group 270:  members (2) 
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/$exit
      -- CP-element group 270: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Sample/ra
      -- 
    ra_2930_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 270_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_0, ack => testConfigure_CP_0_elements(270)); -- 
    -- CP-element group 271:  transition  input  bypass 
    -- CP-element group 271: predecessors 
    -- CP-element group 271: 	61 
    -- CP-element group 271: successors 
    -- CP-element group 271: 	272 
    -- CP-element group 271:  members (2) 
      -- CP-element group 271: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/$exit
      -- CP-element group 271: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/Update/ca
      -- 
    ca_2935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 271_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_267_inst_ack_1, ack => testConfigure_CP_0_elements(271)); -- 
    -- CP-element group 272:  join  transition  output  bypass 
    -- CP-element group 272: predecessors 
    -- CP-element group 272: 	270 
    -- CP-element group 272: 	271 
    -- CP-element group 272: successors 
    -- CP-element group 272: 	273 
    -- CP-element group 272:  members (5) 
      -- CP-element group 272: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_267/SplitProtocol/$exit
      -- CP-element group 272: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- 
    phi_stmt_264_req_2936_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_2936_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(272), ack => phi_stmt_264_req_0); -- 
    testConfigure_cp_element_group_272: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_272"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(270) & testConfigure_CP_0_elements(271);
      gj_testConfigure_cp_element_group_272 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(272), clk => clk, reset => reset); --
    end block;
    -- CP-element group 273:  join  transition  bypass 
    -- CP-element group 273: predecessors 
    -- CP-element group 273: 	269 
    -- CP-element group 273: 	272 
    -- CP-element group 273: successors 
    -- CP-element group 273: 	281 
    -- CP-element group 273:  members (1) 
      -- CP-element group 273: 	 branch_block_stmt_32/bbx_xnph221_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_273: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_273"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(269) & testConfigure_CP_0_elements(272);
      gj_testConfigure_cp_element_group_273 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(273), clk => clk, reset => reset); --
    end block;
    -- CP-element group 274:  transition  input  bypass 
    -- CP-element group 274: predecessors 
    -- CP-element group 274: 	72 
    -- CP-element group 274: successors 
    -- CP-element group 274: 	276 
    -- CP-element group 274:  members (2) 
      -- CP-element group 274: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/$exit
      -- CP-element group 274: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Sample/ra
      -- 
    ra_2956_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 274_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_0, ack => testConfigure_CP_0_elements(274)); -- 
    -- CP-element group 275:  transition  input  bypass 
    -- CP-element group 275: predecessors 
    -- CP-element group 275: 	72 
    -- CP-element group 275: successors 
    -- CP-element group 275: 	276 
    -- CP-element group 275:  members (2) 
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/$exit
      -- CP-element group 275: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/Update/ca
      -- 
    ca_2961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 275_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_263_inst_ack_1, ack => testConfigure_CP_0_elements(275)); -- 
    -- CP-element group 276:  join  transition  output  bypass 
    -- CP-element group 276: predecessors 
    -- CP-element group 276: 	274 
    -- CP-element group 276: 	275 
    -- CP-element group 276: successors 
    -- CP-element group 276: 	280 
    -- CP-element group 276:  members (5) 
      -- CP-element group 276: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_sources/type_cast_263/SplitProtocol/$exit
      -- CP-element group 276: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_257/phi_stmt_257_req
      -- 
    phi_stmt_257_req_2962_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_257_req_2962_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(276), ack => phi_stmt_257_req_1); -- 
    testConfigure_cp_element_group_276: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_276"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(274) & testConfigure_CP_0_elements(275);
      gj_testConfigure_cp_element_group_276 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(276), clk => clk, reset => reset); --
    end block;
    -- CP-element group 277:  transition  input  bypass 
    -- CP-element group 277: predecessors 
    -- CP-element group 277: 	72 
    -- CP-element group 277: successors 
    -- CP-element group 277: 	279 
    -- CP-element group 277:  members (2) 
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/$exit
      -- CP-element group 277: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Sample/ra
      -- 
    ra_2979_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 277_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_0, ack => testConfigure_CP_0_elements(277)); -- 
    -- CP-element group 278:  transition  input  bypass 
    -- CP-element group 278: predecessors 
    -- CP-element group 278: 	72 
    -- CP-element group 278: successors 
    -- CP-element group 278: 	279 
    -- CP-element group 278:  members (2) 
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/$exit
      -- CP-element group 278: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/Update/ca
      -- 
    ca_2984_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 278_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_269_inst_ack_1, ack => testConfigure_CP_0_elements(278)); -- 
    -- CP-element group 279:  join  transition  output  bypass 
    -- CP-element group 279: predecessors 
    -- CP-element group 279: 	277 
    -- CP-element group 279: 	278 
    -- CP-element group 279: successors 
    -- CP-element group 279: 	280 
    -- CP-element group 279:  members (5) 
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_sources/type_cast_269/SplitProtocol/$exit
      -- CP-element group 279: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/phi_stmt_264/phi_stmt_264_req
      -- 
    phi_stmt_264_req_2985_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_264_req_2985_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(279), ack => phi_stmt_264_req_1); -- 
    testConfigure_cp_element_group_279: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_279"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(277) & testConfigure_CP_0_elements(278);
      gj_testConfigure_cp_element_group_279 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(279), clk => clk, reset => reset); --
    end block;
    -- CP-element group 280:  join  transition  bypass 
    -- CP-element group 280: predecessors 
    -- CP-element group 280: 	276 
    -- CP-element group 280: 	279 
    -- CP-element group 280: successors 
    -- CP-element group 280: 	281 
    -- CP-element group 280:  members (1) 
      -- CP-element group 280: 	 branch_block_stmt_32/forx_xbody28_forx_xbody28_PhiReq/$exit
      -- 
    testConfigure_cp_element_group_280: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_280"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(276) & testConfigure_CP_0_elements(279);
      gj_testConfigure_cp_element_group_280 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(280), clk => clk, reset => reset); --
    end block;
    -- CP-element group 281:  merge  fork  transition  place  bypass 
    -- CP-element group 281: predecessors 
    -- CP-element group 281: 	273 
    -- CP-element group 281: 	280 
    -- CP-element group 281: successors 
    -- CP-element group 281: 	282 
    -- CP-element group 281: 	283 
    -- CP-element group 281:  members (2) 
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_256_PhiReqMerge
      -- CP-element group 281: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(281) <= OrReduce(testConfigure_CP_0_elements(273) & testConfigure_CP_0_elements(280));
    -- CP-element group 282:  transition  input  bypass 
    -- CP-element group 282: predecessors 
    -- CP-element group 282: 	281 
    -- CP-element group 282: successors 
    -- CP-element group 282: 	284 
    -- CP-element group 282:  members (1) 
      -- CP-element group 282: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/phi_stmt_257_ack
      -- 
    phi_stmt_257_ack_2990_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 282_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_257_ack_0, ack => testConfigure_CP_0_elements(282)); -- 
    -- CP-element group 283:  transition  input  bypass 
    -- CP-element group 283: predecessors 
    -- CP-element group 283: 	281 
    -- CP-element group 283: successors 
    -- CP-element group 283: 	284 
    -- CP-element group 283:  members (1) 
      -- CP-element group 283: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/phi_stmt_264_ack
      -- 
    phi_stmt_264_ack_2991_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 283_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_264_ack_0, ack => testConfigure_CP_0_elements(283)); -- 
    -- CP-element group 284:  join  fork  transition  place  output  bypass 
    -- CP-element group 284: predecessors 
    -- CP-element group 284: 	282 
    -- CP-element group 284: 	283 
    -- CP-element group 284: successors 
    -- CP-element group 284: 	62 
    -- CP-element group 284: 	63 
    -- CP-element group 284: 	65 
    -- CP-element group 284: 	66 
    -- CP-element group 284: 	69 
    -- CP-element group 284:  members (42) 
      -- CP-element group 284: 	 branch_block_stmt_32/merge_stmt_256__exit__
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298__entry__
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_complete/req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_root_address_calculated
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_offset_calculated
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resized_0
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scaled_0
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_computed_0
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/index_resize_req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_resize_0/index_resize_ack
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/scale_rename_req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_index_scale_0/scale_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_final_index_sum_regn/ack
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/$exit
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/sum_rename_req
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/array_obj_ref_273_base_plus_offset/sum_rename_ack
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/addr_of_274_request/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/ptr_deref_277_Update/word_access_complete/word_0/cr
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_sample_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/RPIPE_ConvTranspose_input_pipe_281_Sample/rr
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_update_start_
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/$entry
      -- CP-element group 284: 	 branch_block_stmt_32/assign_stmt_275_to_assign_stmt_298/type_cast_285_Update/cr
      -- CP-element group 284: 	 branch_block_stmt_32/merge_stmt_256_PhiAck/$exit
      -- 
    req_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_274_final_reg_req_0); -- 
    req_801_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_801_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => addr_of_274_final_reg_req_1); -- 
    cr_851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => ptr_deref_277_store_0_req_1); -- 
    rr_860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => RPIPE_ConvTranspose_input_pipe_281_inst_req_0); -- 
    cr_879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(284), ack => type_cast_285_inst_req_1); -- 
    testConfigure_cp_element_group_284: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_284"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(282) & testConfigure_CP_0_elements(283);
      gj_testConfigure_cp_element_group_284 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(284), clk => clk, reset => reset); --
    end block;
    -- CP-element group 285:  transition  input  bypass 
    -- CP-element group 285: predecessors 
    -- CP-element group 285: 	71 
    -- CP-element group 285: successors 
    -- CP-element group 285: 	287 
    -- CP-element group 285:  members (2) 
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/$exit
      -- CP-element group 285: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Sample/ra
      -- 
    ra_3015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 285_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_0, ack => testConfigure_CP_0_elements(285)); -- 
    -- CP-element group 286:  transition  input  bypass 
    -- CP-element group 286: predecessors 
    -- CP-element group 286: 	71 
    -- CP-element group 286: successors 
    -- CP-element group 286: 	287 
    -- CP-element group 286:  members (2) 
      -- CP-element group 286: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/$exit
      -- CP-element group 286: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/Update/ca
      -- 
    ca_3020_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 286_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_309_inst_ack_1, ack => testConfigure_CP_0_elements(286)); -- 
    -- CP-element group 287:  join  transition  place  output  bypass 
    -- CP-element group 287: predecessors 
    -- CP-element group 287: 	285 
    -- CP-element group 287: 	286 
    -- CP-element group 287: successors 
    -- CP-element group 287: 	288 
    -- CP-element group 287:  members (8) 
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_sources/type_cast_309/SplitProtocol/$exit
      -- CP-element group 287: 	 branch_block_stmt_32/forx_xbody28_forx_xend37_PhiReq/phi_stmt_306/phi_stmt_306_req
      -- CP-element group 287: 	 branch_block_stmt_32/merge_stmt_305_PhiReqMerge
      -- CP-element group 287: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/$entry
      -- 
    phi_stmt_306_req_3021_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_306_req_3021_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(287), ack => phi_stmt_306_req_0); -- 
    testConfigure_cp_element_group_287: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_287"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(285) & testConfigure_CP_0_elements(286);
      gj_testConfigure_cp_element_group_287 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(287), clk => clk, reset => reset); --
    end block;
    -- CP-element group 288:  merge  transition  place  input  bypass 
    -- CP-element group 288: predecessors 
    -- CP-element group 288: 	287 
    -- CP-element group 288: successors 
    -- CP-element group 288: 	73 
    -- CP-element group 288:  members (4) 
      -- CP-element group 288: 	 branch_block_stmt_32/merge_stmt_305__exit__
      -- CP-element group 288: 	 branch_block_stmt_32/assign_stmt_313_to_assign_stmt_499__entry__
      -- CP-element group 288: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/$exit
      -- CP-element group 288: 	 branch_block_stmt_32/merge_stmt_305_PhiAck/phi_stmt_306_ack
      -- 
    phi_stmt_306_ack_3026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 288_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_306_ack_0, ack => testConfigure_CP_0_elements(288)); -- 
    -- CP-element group 289:  merge  branch  transition  place  output  bypass 
    -- CP-element group 289: predecessors 
    -- CP-element group 289: 	120 
    -- CP-element group 289: 	166 
    -- CP-element group 289: successors 
    -- CP-element group 289: 	122 
    -- CP-element group 289: 	123 
    -- CP-element group 289:  members (17) 
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_508__exit__
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520__entry__
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520__exit__
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521__entry__
      -- CP-element group 289: 	 branch_block_stmt_32/assign_stmt_514_to_assign_stmt_520/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_dead_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_eval_test/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_eval_test/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_eval_test/branch_req
      -- CP-element group 289: 	 branch_block_stmt_32/R_cmp124208_522_place
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_if_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/if_stmt_521_else_link/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_508_PhiReqMerge
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/$entry
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/$exit
      -- CP-element group 289: 	 branch_block_stmt_32/merge_stmt_508_PhiAck/dummy
      -- 
    branch_req_1579_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1579_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(289), ack => if_stmt_521_branch_req_0); -- 
    testConfigure_CP_0_elements(289) <= OrReduce(testConfigure_CP_0_elements(120) & testConfigure_CP_0_elements(166));
    -- CP-element group 290:  transition  output  delay-element  bypass 
    -- CP-element group 290: predecessors 
    -- CP-element group 290: 	125 
    -- CP-element group 290: successors 
    -- CP-element group 290: 	294 
    -- CP-element group 290:  members (5) 
      -- CP-element group 290: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$exit
      -- CP-element group 290: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_567_konst_delay_trans
      -- CP-element group 290: 	 branch_block_stmt_32/bbx_xnph215_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_req
      -- 
    phi_stmt_563_req_3072_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_563_req_3072_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(290), ack => phi_stmt_563_req_0); -- 
    -- Element group testConfigure_CP_0_elements(290) is a control-delay.
    cp_element_290_delay: control_delay_element  generic map(name => " 290_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(125), ack => testConfigure_CP_0_elements(290), clk => clk, reset =>reset);
    -- CP-element group 291:  transition  input  bypass 
    -- CP-element group 291: predecessors 
    -- CP-element group 291: 	167 
    -- CP-element group 291: successors 
    -- CP-element group 291: 	293 
    -- CP-element group 291:  members (2) 
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/$exit
      -- CP-element group 291: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Sample/ra
      -- 
    ra_3092_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 291_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_0, ack => testConfigure_CP_0_elements(291)); -- 
    -- CP-element group 292:  transition  input  bypass 
    -- CP-element group 292: predecessors 
    -- CP-element group 292: 	167 
    -- CP-element group 292: successors 
    -- CP-element group 292: 	293 
    -- CP-element group 292:  members (2) 
      -- CP-element group 292: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/$exit
      -- CP-element group 292: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/Update/ca
      -- 
    ca_3097_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 292_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_569_inst_ack_1, ack => testConfigure_CP_0_elements(292)); -- 
    -- CP-element group 293:  join  transition  output  bypass 
    -- CP-element group 293: predecessors 
    -- CP-element group 293: 	291 
    -- CP-element group 293: 	292 
    -- CP-element group 293: successors 
    -- CP-element group 293: 	294 
    -- CP-element group 293:  members (6) 
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_sources/type_cast_569/SplitProtocol/$exit
      -- CP-element group 293: 	 branch_block_stmt_32/forx_xbody67_forx_xbody67_PhiReq/phi_stmt_563/phi_stmt_563_req
      -- 
    phi_stmt_563_req_3098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_563_req_3098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(293), ack => phi_stmt_563_req_1); -- 
    testConfigure_cp_element_group_293: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_293"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(291) & testConfigure_CP_0_elements(292);
      gj_testConfigure_cp_element_group_293 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(293), clk => clk, reset => reset); --
    end block;
    -- CP-element group 294:  merge  transition  place  bypass 
    -- CP-element group 294: predecessors 
    -- CP-element group 294: 	290 
    -- CP-element group 294: 	293 
    -- CP-element group 294: successors 
    -- CP-element group 294: 	295 
    -- CP-element group 294:  members (2) 
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_562_PhiReqMerge
      -- CP-element group 294: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(294) <= OrReduce(testConfigure_CP_0_elements(290) & testConfigure_CP_0_elements(293));
    -- CP-element group 295:  fork  transition  place  input  output  bypass 
    -- CP-element group 295: predecessors 
    -- CP-element group 295: 	294 
    -- CP-element group 295: successors 
    -- CP-element group 295: 	126 
    -- CP-element group 295: 	127 
    -- CP-element group 295: 	129 
    -- CP-element group 295: 	130 
    -- CP-element group 295: 	133 
    -- CP-element group 295: 	137 
    -- CP-element group 295: 	141 
    -- CP-element group 295: 	145 
    -- CP-element group 295: 	149 
    -- CP-element group 295: 	153 
    -- CP-element group 295: 	157 
    -- CP-element group 295: 	161 
    -- CP-element group 295: 	164 
    -- CP-element group 295:  members (56) 
      -- CP-element group 295: 	 branch_block_stmt_32/merge_stmt_562__exit__
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725__entry__
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resized_1
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scaled_1
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_computed_1
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/index_resize_req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_resize_1/index_resize_ack
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/scale_rename_req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_index_scale_1/scale_rename_ack
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_update_start
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Sample/req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/array_obj_ref_575_final_index_sum_regn_Update/req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/addr_of_576_complete/req
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_sample_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/RPIPE_ConvTranspose_input_pipe_579_Sample/rr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_583_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_596_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_614_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_632_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_650_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_668_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_686_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/type_cast_704_Update/cr
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_update_start_
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/$entry
      -- CP-element group 295: 	 branch_block_stmt_32/assign_stmt_577_to_assign_stmt_725/ptr_deref_712_Update/word_access_complete/word_0/cr
      -- CP-element group 295: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/$exit
      -- CP-element group 295: 	 branch_block_stmt_32/merge_stmt_562_PhiAck/phi_stmt_563_ack
      -- 
    phi_stmt_563_ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 295_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_563_ack_0, ack => testConfigure_CP_0_elements(295)); -- 
    req_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_575_index_offset_req_0); -- 
    req_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => array_obj_ref_575_index_offset_req_1); -- 
    req_1655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => addr_of_576_final_reg_req_1); -- 
    rr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => RPIPE_ConvTranspose_input_pipe_579_inst_req_0); -- 
    cr_1683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_583_inst_req_1); -- 
    cr_1711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_596_inst_req_1); -- 
    cr_1739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_614_inst_req_1); -- 
    cr_1767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_632_inst_req_1); -- 
    cr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_650_inst_req_1); -- 
    cr_1823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_668_inst_req_1); -- 
    cr_1851_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1851_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_686_inst_req_1); -- 
    cr_1879_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1879_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => type_cast_704_inst_req_1); -- 
    cr_1929_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1929_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(295), ack => ptr_deref_712_store_0_req_1); -- 
    -- CP-element group 296:  transition  output  delay-element  bypass 
    -- CP-element group 296: predecessors 
    -- CP-element group 296: 	169 
    -- CP-element group 296: successors 
    -- CP-element group 296: 	300 
    -- CP-element group 296:  members (5) 
      -- CP-element group 296: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$exit
      -- CP-element group 296: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_777_konst_delay_trans
      -- CP-element group 296: 	 branch_block_stmt_32/bbx_xnph210_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_req
      -- 
    phi_stmt_773_req_3126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_773_req_3126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(296), ack => phi_stmt_773_req_0); -- 
    -- Element group testConfigure_CP_0_elements(296) is a control-delay.
    cp_element_296_delay: control_delay_element  generic map(name => " 296_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(169), ack => testConfigure_CP_0_elements(296), clk => clk, reset =>reset);
    -- CP-element group 297:  transition  input  bypass 
    -- CP-element group 297: predecessors 
    -- CP-element group 297: 	211 
    -- CP-element group 297: successors 
    -- CP-element group 297: 	299 
    -- CP-element group 297:  members (2) 
      -- CP-element group 297: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/$exit
      -- CP-element group 297: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Sample/ra
      -- 
    ra_3146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 297_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_0, ack => testConfigure_CP_0_elements(297)); -- 
    -- CP-element group 298:  transition  input  bypass 
    -- CP-element group 298: predecessors 
    -- CP-element group 298: 	211 
    -- CP-element group 298: successors 
    -- CP-element group 298: 	299 
    -- CP-element group 298:  members (2) 
      -- CP-element group 298: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/$exit
      -- CP-element group 298: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/Update/ca
      -- 
    ca_3151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 298_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_779_inst_ack_1, ack => testConfigure_CP_0_elements(298)); -- 
    -- CP-element group 299:  join  transition  output  bypass 
    -- CP-element group 299: predecessors 
    -- CP-element group 299: 	297 
    -- CP-element group 299: 	298 
    -- CP-element group 299: successors 
    -- CP-element group 299: 	300 
    -- CP-element group 299:  members (6) 
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_sources/type_cast_779/SplitProtocol/$exit
      -- CP-element group 299: 	 branch_block_stmt_32/forx_xbody126_forx_xbody126_PhiReq/phi_stmt_773/phi_stmt_773_req
      -- 
    phi_stmt_773_req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_773_req_3152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(299), ack => phi_stmt_773_req_1); -- 
    testConfigure_cp_element_group_299: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_299"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(297) & testConfigure_CP_0_elements(298);
      gj_testConfigure_cp_element_group_299 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(299), clk => clk, reset => reset); --
    end block;
    -- CP-element group 300:  merge  transition  place  bypass 
    -- CP-element group 300: predecessors 
    -- CP-element group 300: 	296 
    -- CP-element group 300: 	299 
    -- CP-element group 300: successors 
    -- CP-element group 300: 	301 
    -- CP-element group 300:  members (2) 
      -- CP-element group 300: 	 branch_block_stmt_32/merge_stmt_772_PhiReqMerge
      -- CP-element group 300: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(300) <= OrReduce(testConfigure_CP_0_elements(296) & testConfigure_CP_0_elements(299));
    -- CP-element group 301:  fork  transition  place  input  output  bypass 
    -- CP-element group 301: predecessors 
    -- CP-element group 301: 	300 
    -- CP-element group 301: successors 
    -- CP-element group 301: 	170 
    -- CP-element group 301: 	171 
    -- CP-element group 301: 	173 
    -- CP-element group 301: 	174 
    -- CP-element group 301: 	177 
    -- CP-element group 301: 	181 
    -- CP-element group 301: 	185 
    -- CP-element group 301: 	189 
    -- CP-element group 301: 	193 
    -- CP-element group 301: 	197 
    -- CP-element group 301: 	201 
    -- CP-element group 301: 	205 
    -- CP-element group 301: 	208 
    -- CP-element group 301:  members (56) 
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/merge_stmt_772__exit__
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935__entry__
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_878_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/word_0/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_896_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/word_access_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/ptr_deref_922_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_914_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_860_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resized_1
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scaled_1
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_computed_1
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/index_resize_req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_resize_1/index_resize_ack
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/scale_rename_req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_index_scale_1/scale_rename_ack
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_update_start
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Sample/req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/array_obj_ref_785_final_index_sum_regn_Update/req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/addr_of_786_complete/req
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_sample_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/RPIPE_ConvTranspose_input_pipe_789_Sample/rr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_793_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_806_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/$entry
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_824_Update/cr
      -- CP-element group 301: 	 branch_block_stmt_32/assign_stmt_787_to_assign_stmt_935/type_cast_842_update_start_
      -- CP-element group 301: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/$exit
      -- CP-element group 301: 	 branch_block_stmt_32/merge_stmt_772_PhiAck/phi_stmt_773_ack
      -- 
    phi_stmt_773_ack_3157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 301_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_773_ack_0, ack => testConfigure_CP_0_elements(301)); -- 
    cr_2210_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2210_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_896_inst_req_1); -- 
    cr_2182_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2182_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_878_inst_req_1); -- 
    cr_2238_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2238_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_914_inst_req_1); -- 
    cr_2154_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2154_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_860_inst_req_1); -- 
    cr_2288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => ptr_deref_922_store_0_req_1); -- 
    cr_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_842_inst_req_1); -- 
    req_1994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_785_index_offset_req_0); -- 
    req_1999_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1999_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => array_obj_ref_785_index_offset_req_1); -- 
    req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => addr_of_786_final_reg_req_1); -- 
    rr_2023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => RPIPE_ConvTranspose_input_pipe_789_inst_req_0); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2042_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_793_inst_req_1); -- 
    cr_2070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_806_inst_req_1); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(301), ack => type_cast_824_inst_req_1); -- 
    -- CP-element group 302:  merge  place  bypass 
    -- CP-element group 302: predecessors 
    -- CP-element group 302: 	122 
    -- CP-element group 302: 	210 
    -- CP-element group 302: successors 
    -- CP-element group 302: 	303 
    -- CP-element group 302:  members (1) 
      -- CP-element group 302: 	 branch_block_stmt_32/merge_stmt_944_PhiReqMerge
      -- 
    testConfigure_CP_0_elements(302) <= OrReduce(testConfigure_CP_0_elements(122) & testConfigure_CP_0_elements(210));
    -- CP-element group 303:  join  fork  transition  place  output  bypass 
    -- CP-element group 303: predecessors 
    -- CP-element group 303: 	302 
    -- CP-element group 303: successors 
    -- CP-element group 303: 	212 
    -- CP-element group 303: 	213 
    -- CP-element group 303: 	214 
    -- CP-element group 303: 	215 
    -- CP-element group 303: 	216 
    -- CP-element group 303: 	217 
    -- CP-element group 303:  members (84) 
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_32/merge_stmt_944__exit__
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996__entry__
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_word_addrgen/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_word_addrgen/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_plus_offset/sum_rename_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_plus_offset/sum_rename_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_plus_offset/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_plus_offset/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_addr_resize/base_resize_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_addr_resize/base_resize_req
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_addr_resize/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_addr_resize/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_address_resized
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_root_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_word_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_base_address_calculated
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_update_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_979_sample_start_
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/word_access_complete/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Update/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/word_0/rr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/word_access_start/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/word_0/cr
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_955_Update/word_access_complete/word_0/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_Sample/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_word_addrgen/root_register_ack
      -- CP-element group 303: 	 branch_block_stmt_32/assign_stmt_952_to_assign_stmt_996/ptr_deref_967_word_addrgen/root_register_req
      -- CP-element group 303: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/$entry
      -- CP-element group 303: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/$exit
      -- CP-element group 303: 	 branch_block_stmt_32/merge_stmt_944_PhiAck/dummy
      -- 
    cr_2455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_979_load_0_req_1); -- 
    rr_2344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_955_load_0_req_0); -- 
    rr_2444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_979_load_0_req_0); -- 
    cr_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_967_load_0_req_1); -- 
    rr_2394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_967_load_0_req_0); -- 
    cr_2355_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2355_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(303), ack => ptr_deref_955_load_0_req_1); -- 
    testConfigure_CP_0_elements(303) <= testConfigure_CP_0_elements(302);
    -- CP-element group 304:  transition  output  delay-element  bypass 
    -- CP-element group 304: predecessors 
    -- CP-element group 304: 	222 
    -- CP-element group 304: successors 
    -- CP-element group 304: 	308 
    -- CP-element group 304:  members (5) 
      -- CP-element group 304: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$exit
      -- CP-element group 304: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1045_konst_delay_trans
      -- CP-element group 304: 	 branch_block_stmt_32/bbx_xnph_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_req
      -- 
    phi_stmt_1041_req_3203_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1041_req_3203_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(304), ack => phi_stmt_1041_req_0); -- 
    -- Element group testConfigure_CP_0_elements(304) is a control-delay.
    cp_element_304_delay: control_delay_element  generic map(name => " 304_delay", delay_value => 1)  port map(req => testConfigure_CP_0_elements(222), ack => testConfigure_CP_0_elements(304), clk => clk, reset =>reset);
    -- CP-element group 305:  transition  input  bypass 
    -- CP-element group 305: predecessors 
    -- CP-element group 305: 	231 
    -- CP-element group 305: successors 
    -- CP-element group 305: 	307 
    -- CP-element group 305:  members (2) 
      -- CP-element group 305: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Sample/$exit
      -- CP-element group 305: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Sample/ra
      -- 
    ra_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 305_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1047_inst_ack_0, ack => testConfigure_CP_0_elements(305)); -- 
    -- CP-element group 306:  transition  input  bypass 
    -- CP-element group 306: predecessors 
    -- CP-element group 306: 	231 
    -- CP-element group 306: successors 
    -- CP-element group 306: 	307 
    -- CP-element group 306:  members (2) 
      -- CP-element group 306: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Update/$exit
      -- CP-element group 306: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/Update/ca
      -- 
    ca_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 306_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1047_inst_ack_1, ack => testConfigure_CP_0_elements(306)); -- 
    -- CP-element group 307:  join  transition  output  bypass 
    -- CP-element group 307: predecessors 
    -- CP-element group 307: 	305 
    -- CP-element group 307: 	306 
    -- CP-element group 307: successors 
    -- CP-element group 307: 	308 
    -- CP-element group 307:  members (6) 
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_sources/type_cast_1047/SplitProtocol/$exit
      -- CP-element group 307: 	 branch_block_stmt_32/forx_xbody193_forx_xbody193_PhiReq/phi_stmt_1041/phi_stmt_1041_req
      -- 
    phi_stmt_1041_req_3229_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1041_req_3229_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(307), ack => phi_stmt_1041_req_1); -- 
    testConfigure_cp_element_group_307: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "testConfigure_cp_element_group_307"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= testConfigure_CP_0_elements(305) & testConfigure_CP_0_elements(306);
      gj_testConfigure_cp_element_group_307 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => testConfigure_CP_0_elements(307), clk => clk, reset => reset); --
    end block;
    -- CP-element group 308:  merge  transition  place  bypass 
    -- CP-element group 308: predecessors 
    -- CP-element group 308: 	304 
    -- CP-element group 308: 	307 
    -- CP-element group 308: successors 
    -- CP-element group 308: 	309 
    -- CP-element group 308:  members (2) 
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1040_PhiReqMerge
      -- CP-element group 308: 	 branch_block_stmt_32/merge_stmt_1040_PhiAck/$entry
      -- 
    testConfigure_CP_0_elements(308) <= OrReduce(testConfigure_CP_0_elements(304) & testConfigure_CP_0_elements(307));
    -- CP-element group 309:  fork  transition  place  input  output  bypass 
    -- CP-element group 309: predecessors 
    -- CP-element group 309: 	308 
    -- CP-element group 309: successors 
    -- CP-element group 309: 	223 
    -- CP-element group 309: 	224 
    -- CP-element group 309: 	226 
    -- CP-element group 309: 	228 
    -- CP-element group 309:  members (29) 
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_complete/req
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/merge_stmt_1040__exit__
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071__entry__
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Update/req
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_resized_1
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Sample/req
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_Sample/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/addr_of_1054_update_start_
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_final_index_sum_regn_update_start
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_scale_1/scale_rename_ack
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_scale_1/scale_rename_req
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_scale_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_scale_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_resize_1/index_resize_ack
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/word_0/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_resize_1/$entry
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_computed_1
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_resize_1/index_resize_req
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_resize_1/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/array_obj_ref_1053_index_scaled_1
      -- CP-element group 309: 	 branch_block_stmt_32/assign_stmt_1055_to_assign_stmt_1071/ptr_deref_1057_Update/word_access_complete/word_0/cr
      -- CP-element group 309: 	 branch_block_stmt_32/merge_stmt_1040_PhiAck/$exit
      -- CP-element group 309: 	 branch_block_stmt_32/merge_stmt_1040_PhiAck/phi_stmt_1041_ack
      -- 
    phi_stmt_1041_ack_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 309_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1041_ack_0, ack => testConfigure_CP_0_elements(309)); -- 
    req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2545_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => addr_of_1054_final_reg_req_1); -- 
    req_2530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1053_index_offset_req_1); -- 
    req_2525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => array_obj_ref_1053_index_offset_req_0); -- 
    cr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2595_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(309), ack => ptr_deref_1057_store_0_req_1); -- 
    -- CP-element group 310:  merge  fork  transition  place  output  bypass 
    -- CP-element group 310: predecessors 
    -- CP-element group 310: 	220 
    -- CP-element group 310: 	230 
    -- CP-element group 310: successors 
    -- CP-element group 310: 	232 
    -- CP-element group 310: 	233 
    -- CP-element group 310:  members (13) 
      -- CP-element group 310: 	 branch_block_stmt_32/merge_stmt_1080__exit__
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084__entry__
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_sample_start_
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_update_start_
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Sample/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Sample/rr
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Update/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/assign_stmt_1084/type_cast_1083_Update/cr
      -- CP-element group 310: 	 branch_block_stmt_32/merge_stmt_1080_PhiReqMerge
      -- CP-element group 310: 	 branch_block_stmt_32/merge_stmt_1080_PhiAck/$entry
      -- CP-element group 310: 	 branch_block_stmt_32/merge_stmt_1080_PhiAck/$exit
      -- CP-element group 310: 	 branch_block_stmt_32/merge_stmt_1080_PhiAck/dummy
      -- 
    rr_2626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1083_inst_req_0); -- 
    cr_2631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => testConfigure_CP_0_elements(310), ack => type_cast_1083_inst_req_1); -- 
    testConfigure_CP_0_elements(310) <= OrReduce(testConfigure_CP_0_elements(220) & testConfigure_CP_0_elements(230));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_indvar240_784_resized : std_logic_vector(10 downto 0);
    signal R_indvar240_784_scaled : std_logic_vector(10 downto 0);
    signal R_indvar250_574_resized : std_logic_vector(13 downto 0);
    signal R_indvar250_574_scaled : std_logic_vector(13 downto 0);
    signal R_indvar260_272_resized : std_logic_vector(0 downto 0);
    signal R_indvar260_272_scaled : std_logic_vector(0 downto 0);
    signal R_indvar263_203_resized : std_logic_vector(6 downto 0);
    signal R_indvar263_203_scaled : std_logic_vector(6 downto 0);
    signal R_indvar268_100_resized : std_logic_vector(6 downto 0);
    signal R_indvar268_100_scaled : std_logic_vector(6 downto 0);
    signal R_indvar_1052_resized : std_logic_vector(13 downto 0);
    signal R_indvar_1052_scaled : std_logic_vector(13 downto 0);
    signal STORE_padding_311_data_0 : std_logic_vector(15 downto 0);
    signal STORE_padding_311_word_address_0 : std_logic_vector(0 downto 0);
    signal add104_692 : std_logic_vector(63 downto 0);
    signal add110_710 : std_logic_vector(63 downto 0);
    signal add136_812 : std_logic_vector(63 downto 0);
    signal add142_830 : std_logic_vector(63 downto 0);
    signal add148_848 : std_logic_vector(63 downto 0);
    signal add154_866 : std_logic_vector(63 downto 0);
    signal add160_884 : std_logic_vector(63 downto 0);
    signal add166_902 : std_logic_vector(63 downto 0);
    signal add172_920 : std_logic_vector(63 downto 0);
    signal add80_620 : std_logic_vector(63 downto 0);
    signal add86_638 : std_logic_vector(63 downto 0);
    signal add92_656 : std_logic_vector(63 downto 0);
    signal add98_674 : std_logic_vector(63 downto 0);
    signal add_602 : std_logic_vector(63 downto 0);
    signal array_obj_ref_101_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_101_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1053_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1053_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1053_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1053_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1053_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1053_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_204_constant_part_of_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_offset_scale_factor_1 : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_204_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_273_final_offset : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_offset_scale_factor_0 : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_resized_base_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_273_root_address : std_logic_vector(0 downto 0);
    signal array_obj_ref_575_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_575_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_785_constant_part_of_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_offset_scale_factor_1 : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_785_root_address : std_logic_vector(10 downto 0);
    signal arrayidx114_577 : std_logic_vector(31 downto 0);
    signal arrayidx176_787 : std_logic_vector(31 downto 0);
    signal arrayidx196_1055 : std_logic_vector(31 downto 0);
    signal arrayidx19_206 : std_logic_vector(31 downto 0);
    signal arrayidx33_275 : std_logic_vector(31 downto 0);
    signal arrayidx_103 : std_logic_vector(31 downto 0);
    signal call101_683 : std_logic_vector(7 downto 0);
    signal call107_701 : std_logic_vector(7 downto 0);
    signal call129_790 : std_logic_vector(7 downto 0);
    signal call133_803 : std_logic_vector(7 downto 0);
    signal call139_821 : std_logic_vector(7 downto 0);
    signal call145_839 : std_logic_vector(7 downto 0);
    signal call151_857 : std_logic_vector(7 downto 0);
    signal call157_875 : std_logic_vector(7 downto 0);
    signal call15_209 : std_logic_vector(7 downto 0);
    signal call163_893 : std_logic_vector(7 downto 0);
    signal call169_911 : std_logic_vector(7 downto 0);
    signal call29217_250 : std_logic_vector(7 downto 0);
    signal call29_282 : std_logic_vector(7 downto 0);
    signal call3228_59 : std_logic_vector(7 downto 0);
    signal call3_131 : std_logic_vector(7 downto 0);
    signal call40_316 : std_logic_vector(7 downto 0);
    signal call42_335 : std_logic_vector(7 downto 0);
    signal call44_354 : std_logic_vector(7 downto 0);
    signal call69_580 : std_logic_vector(7 downto 0);
    signal call72_593 : std_logic_vector(7 downto 0);
    signal call77_611 : std_logic_vector(7 downto 0);
    signal call83_629 : std_logic_vector(7 downto 0);
    signal call89_647 : std_logic_vector(7 downto 0);
    signal call95_665 : std_logic_vector(7 downto 0);
    signal call_35 : std_logic_vector(7 downto 0);
    signal cmp12223_172 : std_logic_vector(0 downto 0);
    signal cmp124208_520 : std_logic_vector(0 downto 0);
    signal cmp12_238 : std_logic_vector(0 downto 0);
    signal cmp191204_996 : std_logic_vector(0 downto 0);
    signal cmp227_56 : std_logic_vector(0 downto 0);
    signal cmp65213_499 : std_logic_vector(0 downto 0);
    signal cmp_128 : std_logic_vector(0 downto 0);
    signal conv103_687 : std_logic_vector(63 downto 0);
    signal conv109_705 : std_logic_vector(63 downto 0);
    signal conv130_794 : std_logic_vector(63 downto 0);
    signal conv135_807 : std_logic_vector(63 downto 0);
    signal conv141_825 : std_logic_vector(63 downto 0);
    signal conv147_843 : std_logic_vector(63 downto 0);
    signal conv153_861 : std_logic_vector(63 downto 0);
    signal conv159_879 : std_logic_vector(63 downto 0);
    signal conv165_897 : std_logic_vector(63 downto 0);
    signal conv16_213 : std_logic_vector(31 downto 0);
    signal conv171_915 : std_logic_vector(63 downto 0);
    signal conv30218_254 : std_logic_vector(15 downto 0);
    signal conv30220_264 : std_logic_vector(15 downto 0);
    signal conv30_286 : std_logic_vector(15 downto 0);
    signal conv30x_xlcssa_306 : std_logic_vector(15 downto 0);
    signal conv41_320 : std_logic_vector(31 downto 0);
    signal conv4229_63 : std_logic_vector(31 downto 0);
    signal conv4231_80 : std_logic_vector(31 downto 0);
    signal conv43_339 : std_logic_vector(31 downto 0);
    signal conv45_358 : std_logic_vector(31 downto 0);
    signal conv4_135 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa1_143 : std_logic_vector(31 downto 0);
    signal conv4x_xlcssa_150 : std_logic_vector(31 downto 0);
    signal conv51_420 : std_logic_vector(63 downto 0);
    signal conv60_487 : std_logic_vector(63 downto 0);
    signal conv70_584 : std_logic_vector(63 downto 0);
    signal conv74_597 : std_logic_vector(63 downto 0);
    signal conv79_615 : std_logic_vector(63 downto 0);
    signal conv85_633 : std_logic_vector(63 downto 0);
    signal conv91_651 : std_logic_vector(63 downto 0);
    signal conv97_669 : std_logic_vector(63 downto 0);
    signal conv_39 : std_logic_vector(31 downto 0);
    signal exitcond10_725 : std_logic_vector(0 downto 0);
    signal exitcond19_935 : std_logic_vector(0 downto 0);
    signal exitcond20_1071 : std_logic_vector(0 downto 0);
    signal exitcond_298 : std_logic_vector(0 downto 0);
    signal iNsTr_13_119 : std_logic_vector(31 downto 0);
    signal iNsTr_1_45 : std_logic_vector(31 downto 0);
    signal iNsTr_21_229 : std_logic_vector(31 downto 0);
    signal iNsTr_26_328 : std_logic_vector(31 downto 0);
    signal iNsTr_29_347 : std_logic_vector(31 downto 0);
    signal iNsTr_32_366 : std_logic_vector(31 downto 0);
    signal iNsTr_34_378 : std_logic_vector(31 downto 0);
    signal iNsTr_35_390 : std_logic_vector(31 downto 0);
    signal iNsTr_36_402 : std_logic_vector(31 downto 0);
    signal iNsTr_37_428 : std_logic_vector(31 downto 0);
    signal iNsTr_38_440 : std_logic_vector(31 downto 0);
    signal iNsTr_39_452 : std_logic_vector(31 downto 0);
    signal iNsTr_40_464 : std_logic_vector(31 downto 0);
    signal iNsTr_45_952 : std_logic_vector(31 downto 0);
    signal iNsTr_46_964 : std_logic_vector(31 downto 0);
    signal iNsTr_47_976 : std_logic_vector(31 downto 0);
    signal iNsTr_5_162 : std_logic_vector(31 downto 0);
    signal iNsTr_60_1025 : std_logic_vector(63 downto 0);
    signal inc22_199 : std_logic_vector(31 downto 0);
    signal inc_96 : std_logic_vector(31 downto 0);
    signal indvar240_773 : std_logic_vector(63 downto 0);
    signal indvar250_563 : std_logic_vector(63 downto 0);
    signal indvar260_257 : std_logic_vector(63 downto 0);
    signal indvar263_182 : std_logic_vector(63 downto 0);
    signal indvar268_73 : std_logic_vector(63 downto 0);
    signal indvar_1041 : std_logic_vector(63 downto 0);
    signal indvarx_xnext241_930 : std_logic_vector(63 downto 0);
    signal indvarx_xnext251_720 : std_logic_vector(63 downto 0);
    signal indvarx_xnext261_292 : std_logic_vector(63 downto 0);
    signal indvarx_xnext_1066 : std_logic_vector(63 downto 0);
    signal mul184_985 : std_logic_vector(31 downto 0);
    signal mul186_990 : std_logic_vector(31 downto 0);
    signal mul50_416 : std_logic_vector(31 downto 0);
    signal mul55_473 : std_logic_vector(31 downto 0);
    signal mul57_478 : std_logic_vector(31 downto 0);
    signal mul59_483 : std_logic_vector(31 downto 0);
    signal mul_411 : std_logic_vector(31 downto 0);
    signal ptr_deref_1057_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_1057_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1057_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1057_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_1057_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1057_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_105_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_105_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_105_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_105_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_105_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_122_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_122_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_164_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_164_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_164_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_164_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_164_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_164_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_215_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_215_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_215_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_215_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_215_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_215_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_232_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_232_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_232_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_232_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_232_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_277_data_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_277_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_277_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_277_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_277_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_277_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_330_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_330_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_330_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_330_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_330_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_330_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_349_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_349_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_349_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_349_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_349_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_349_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_368_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_368_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_368_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_368_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_368_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_368_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_381_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_381_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_393_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_393_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_393_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_393_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_393_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_405_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_405_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_405_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_405_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_405_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_431_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_431_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_431_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_431_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_431_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_443_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_443_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_443_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_443_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_443_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_455_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_455_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_455_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_455_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_455_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_467_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_467_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_467_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_467_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_467_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_47_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_47_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_47_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_47_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_712_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_712_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_712_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_712_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_712_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_712_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_922_data_0 : std_logic_vector(63 downto 0);
    signal ptr_deref_922_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_922_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_922_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_922_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_922_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_955_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_955_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_955_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_955_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_955_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_967_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_967_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_967_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_967_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_967_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_979_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_979_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_979_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_979_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_979_word_offset_0 : std_logic_vector(6 downto 0);
    signal shl100_680 : std_logic_vector(63 downto 0);
    signal shl106_698 : std_logic_vector(63 downto 0);
    signal shl132_800 : std_logic_vector(63 downto 0);
    signal shl138_818 : std_logic_vector(63 downto 0);
    signal shl144_836 : std_logic_vector(63 downto 0);
    signal shl150_854 : std_logic_vector(63 downto 0);
    signal shl156_872 : std_logic_vector(63 downto 0);
    signal shl162_890 : std_logic_vector(63 downto 0);
    signal shl168_908 : std_logic_vector(63 downto 0);
    signal shl76_608 : std_logic_vector(63 downto 0);
    signal shl82_626 : std_logic_vector(63 downto 0);
    signal shl88_644 : std_logic_vector(63 downto 0);
    signal shl94_662 : std_logic_vector(63 downto 0);
    signal shl_590 : std_logic_vector(63 downto 0);
    signal shr123207x_xmask_514 : std_logic_vector(63 downto 0);
    signal shr212x_xmask_493 : std_logic_vector(63 downto 0);
    signal tmp11_233 : std_logic_vector(31 downto 0);
    signal tmp12_737 : std_logic_vector(31 downto 0);
    signal tmp13_742 : std_logic_vector(31 downto 0);
    signal tmp14_747 : std_logic_vector(31 downto 0);
    signal tmp15_751 : std_logic_vector(63 downto 0);
    signal tmp16_757 : std_logic_vector(63 downto 0);
    signal tmp17_763 : std_logic_vector(0 downto 0);
    signal tmp182_956 : std_logic_vector(31 downto 0);
    signal tmp183_968 : std_logic_vector(31 downto 0);
    signal tmp185_980 : std_logic_vector(31 downto 0);
    signal tmp1_123 : std_logic_vector(31 downto 0);
    signal tmp235_1009 : std_logic_vector(31 downto 0);
    signal tmp235x_xop_1021 : std_logic_vector(31 downto 0);
    signal tmp236_1015 : std_logic_vector(0 downto 0);
    signal tmp239_1038 : std_logic_vector(63 downto 0);
    signal tmp265_223 : std_logic_vector(63 downto 0);
    signal tmp270_113 : std_logic_vector(63 downto 0);
    signal tmp3_195 : std_logic_vector(63 downto 0);
    signal tmp47_382 : std_logic_vector(31 downto 0);
    signal tmp48_394 : std_logic_vector(31 downto 0);
    signal tmp49_406 : std_logic_vector(31 downto 0);
    signal tmp53_432 : std_logic_vector(31 downto 0);
    signal tmp54_444 : std_logic_vector(31 downto 0);
    signal tmp56_456 : std_logic_vector(31 downto 0);
    signal tmp58_468 : std_logic_vector(31 downto 0);
    signal tmp5_532 : std_logic_vector(31 downto 0);
    signal tmp6_537 : std_logic_vector(31 downto 0);
    signal tmp7_541 : std_logic_vector(63 downto 0);
    signal tmp8_547 : std_logic_vector(63 downto 0);
    signal tmp9_553 : std_logic_vector(0 downto 0);
    signal tmp_92 : std_logic_vector(63 downto 0);
    signal type_cast_1007_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1013_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1019_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1029_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1036_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1045_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1047_wire : std_logic_vector(63 downto 0);
    signal type_cast_1059_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1064_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_111_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_146_wire : std_logic_vector(31 downto 0);
    signal type_cast_153_wire : std_logic_vector(31 downto 0);
    signal type_cast_155_wire : std_logic_vector(31 downto 0);
    signal type_cast_170_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_185_wire : std_logic_vector(63 downto 0);
    signal type_cast_188_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_193_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_221_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_261_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_263_wire : std_logic_vector(63 downto 0);
    signal type_cast_267_wire : std_logic_vector(15 downto 0);
    signal type_cast_269_wire : std_logic_vector(15 downto 0);
    signal type_cast_290_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_296_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_309_wire : std_logic_vector(15 downto 0);
    signal type_cast_491_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_497_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_512_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_518_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_53_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_545_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_551_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_558_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_567_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_569_wire : std_logic_vector(63 downto 0);
    signal type_cast_588_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_606_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_624_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_642_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_660_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_718_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_761_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_76_wire : std_logic_vector(63 downto 0);
    signal type_cast_777_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_779_wire : std_logic_vector(63 downto 0);
    signal type_cast_798_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_79_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_816_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_834_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_83_wire : std_logic_vector(31 downto 0);
    signal type_cast_852_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_85_wire : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_888_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_90_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_928_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_994_wire_constant : std_logic_vector(31 downto 0);
    signal umax18_770 : std_logic_vector(63 downto 0);
    signal umax_560 : std_logic_vector(63 downto 0);
    signal xx_xop_1031 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    STORE_padding_311_word_address_0 <= "0";
    array_obj_ref_101_constant_part_of_offset <= "0000010";
    array_obj_ref_101_offset_scale_factor_0 <= "1000000";
    array_obj_ref_101_offset_scale_factor_1 <= "0000001";
    array_obj_ref_101_resized_base_address <= "0000000";
    array_obj_ref_1053_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1053_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_1053_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1053_resized_base_address <= "00000000000000";
    array_obj_ref_204_constant_part_of_offset <= "0000010";
    array_obj_ref_204_offset_scale_factor_0 <= "1000000";
    array_obj_ref_204_offset_scale_factor_1 <= "0000001";
    array_obj_ref_204_resized_base_address <= "0000000";
    array_obj_ref_273_offset_scale_factor_0 <= "1";
    array_obj_ref_273_resized_base_address <= "0";
    array_obj_ref_575_constant_part_of_offset <= "00000000000000";
    array_obj_ref_575_offset_scale_factor_0 <= "00000000000000";
    array_obj_ref_575_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_575_resized_base_address <= "00000000000000";
    array_obj_ref_785_constant_part_of_offset <= "00000100001";
    array_obj_ref_785_offset_scale_factor_0 <= "10000000000";
    array_obj_ref_785_offset_scale_factor_1 <= "00000000001";
    array_obj_ref_785_resized_base_address <= "00000000000";
    iNsTr_13_119 <= "00000000000000000000000000000001";
    iNsTr_1_45 <= "00000000000000000000000000000001";
    iNsTr_21_229 <= "00000000000000000000000000000001";
    iNsTr_26_328 <= "00000000000000000000000000000010";
    iNsTr_29_347 <= "00000000000000000000000000000011";
    iNsTr_32_366 <= "00000000000000000000000000000100";
    iNsTr_34_378 <= "00000000000000000000000000000010";
    iNsTr_35_390 <= "00000000000000000000000000000011";
    iNsTr_36_402 <= "00000000000000000000000000000100";
    iNsTr_37_428 <= "00000000000000000000000000000010";
    iNsTr_38_440 <= "00000000000000000000000000000011";
    iNsTr_39_452 <= "00000000000000000000000000000100";
    iNsTr_40_464 <= "00000000000000000000000000000101";
    iNsTr_45_952 <= "00000000000000000000000000000010";
    iNsTr_46_964 <= "00000000000000000000000000000011";
    iNsTr_47_976 <= "00000000000000000000000000000100";
    iNsTr_5_162 <= "00000000000000000000000000000001";
    ptr_deref_1057_word_offset_0 <= "00000000000000";
    ptr_deref_105_word_offset_0 <= "0000000";
    ptr_deref_122_word_offset_0 <= "0000000";
    ptr_deref_164_word_offset_0 <= "0000000";
    ptr_deref_215_word_offset_0 <= "0000000";
    ptr_deref_232_word_offset_0 <= "0000000";
    ptr_deref_277_word_offset_0 <= "0";
    ptr_deref_330_word_offset_0 <= "0000000";
    ptr_deref_349_word_offset_0 <= "0000000";
    ptr_deref_368_word_offset_0 <= "0000000";
    ptr_deref_381_word_offset_0 <= "0000000";
    ptr_deref_393_word_offset_0 <= "0000000";
    ptr_deref_405_word_offset_0 <= "0000000";
    ptr_deref_431_word_offset_0 <= "0000000";
    ptr_deref_443_word_offset_0 <= "0000000";
    ptr_deref_455_word_offset_0 <= "0000000";
    ptr_deref_467_word_offset_0 <= "0000000";
    ptr_deref_47_word_offset_0 <= "0000000";
    ptr_deref_712_word_offset_0 <= "00000000000000";
    ptr_deref_922_word_offset_0 <= "00000000000";
    ptr_deref_955_word_offset_0 <= "0000000";
    ptr_deref_967_word_offset_0 <= "0000000";
    ptr_deref_979_word_offset_0 <= "0000000";
    type_cast_1007_wire_constant <= "00000000000000000000000000000010";
    type_cast_1013_wire_constant <= "00000000000000000000000000000001";
    type_cast_1019_wire_constant <= "11111111111111111111111111111111";
    type_cast_1029_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1036_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1045_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1059_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1064_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_111_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_170_wire_constant <= "00000000000000000000000000000000";
    type_cast_188_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_193_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_221_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_261_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_290_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_296_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_491_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_497_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_512_wire_constant <= "0000000000000000000000000000000011111111111111111111111111111100";
    type_cast_518_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_53_wire_constant <= "00000000";
    type_cast_545_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_551_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_558_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_567_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_588_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_606_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_624_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_642_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_660_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_718_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_755_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000010";
    type_cast_761_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_777_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_798_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_79_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_816_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_834_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_852_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_870_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_888_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_906_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_90_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_928_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_994_wire_constant <= "00000000000000000000000000000011";
    phi_stmt_1041: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1045_wire_constant & type_cast_1047_wire;
      req <= phi_stmt_1041_req_0 & phi_stmt_1041_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1041",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1041_ack_0,
          idata => idata,
          odata => indvar_1041,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1041
    phi_stmt_143: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_146_wire;
      req(0) <= phi_stmt_143_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_143",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_143_ack_0,
          idata => idata,
          odata => conv4x_xlcssa1_143,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_143
    phi_stmt_150: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_153_wire & type_cast_155_wire;
      req <= phi_stmt_150_req_0 & phi_stmt_150_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_150",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_150_ack_0,
          idata => idata,
          odata => conv4x_xlcssa_150,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_150
    phi_stmt_182: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_185_wire & type_cast_188_wire_constant;
      req <= phi_stmt_182_req_0 & phi_stmt_182_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_182",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_182_ack_0,
          idata => idata,
          odata => indvar263_182,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_182
    phi_stmt_257: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_261_wire_constant & type_cast_263_wire;
      req <= phi_stmt_257_req_0 & phi_stmt_257_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_257",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_257_ack_0,
          idata => idata,
          odata => indvar260_257,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_257
    phi_stmt_264: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_267_wire & type_cast_269_wire;
      req <= phi_stmt_264_req_0 & phi_stmt_264_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_264",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_264_ack_0,
          idata => idata,
          odata => conv30220_264,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_264
    phi_stmt_306: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_309_wire;
      req(0) <= phi_stmt_306_req_0;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_306",
          num_reqs => 1,
          bypass_flag => false,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_306_ack_0,
          idata => idata,
          odata => conv30x_xlcssa_306,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_306
    phi_stmt_563: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_567_wire_constant & type_cast_569_wire;
      req <= phi_stmt_563_req_0 & phi_stmt_563_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_563",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_563_ack_0,
          idata => idata,
          odata => indvar250_563,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_563
    phi_stmt_73: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_76_wire & type_cast_79_wire_constant;
      req <= phi_stmt_73_req_0 & phi_stmt_73_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_73",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_73_ack_0,
          idata => idata,
          odata => indvar268_73,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_73
    phi_stmt_773: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_777_wire_constant & type_cast_779_wire;
      req <= phi_stmt_773_req_0 & phi_stmt_773_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_773",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_773_ack_0,
          idata => idata,
          odata => indvar240_773,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_773
    phi_stmt_80: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_83_wire & type_cast_85_wire;
      req <= phi_stmt_80_req_0 & phi_stmt_80_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_80",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_80_ack_0,
          idata => idata,
          odata => conv4231_80,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_80
    -- flow-through select operator MUX_1037_inst
    tmp239_1038 <= xx_xop_1031 when (tmp236_1015(0) /=  '0') else type_cast_1036_wire_constant;
    -- flow-through select operator MUX_559_inst
    umax_560 <= tmp8_547 when (tmp9_553(0) /=  '0') else type_cast_558_wire_constant;
    -- flow-through select operator MUX_769_inst
    umax18_770 <= tmp16_757 when (tmp17_763(0) /=  '0') else type_cast_768_wire_constant;
    addr_of_102_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_102_final_reg_req_0;
      addr_of_102_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_102_final_reg_req_1;
      addr_of_102_final_reg_ack_1<= rack(0);
      addr_of_102_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_102_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_101_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx_103,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_1054_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_1054_final_reg_req_0;
      addr_of_1054_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_1054_final_reg_req_1;
      addr_of_1054_final_reg_ack_1<= rack(0);
      addr_of_1054_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_1054_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_1053_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx196_1055,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_205_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_205_final_reg_req_0;
      addr_of_205_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_205_final_reg_req_1;
      addr_of_205_final_reg_ack_1<= rack(0);
      addr_of_205_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_205_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_204_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx19_206,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_274_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_274_final_reg_req_0;
      addr_of_274_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_274_final_reg_req_1;
      addr_of_274_final_reg_ack_1<= rack(0);
      addr_of_274_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_274_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_273_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx33_275,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_576_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_576_final_reg_req_0;
      addr_of_576_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_576_final_reg_req_1;
      addr_of_576_final_reg_ack_1<= rack(0);
      addr_of_576_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_576_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 14,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_575_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx114_577,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    addr_of_786_final_reg_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= addr_of_786_final_reg_req_0;
      addr_of_786_final_reg_ack_0<= wack(0);
      rreq(0) <= addr_of_786_final_reg_req_1;
      addr_of_786_final_reg_ack_1<= rack(0);
      addr_of_786_final_reg : InterlockBuffer generic map ( -- 
        name => "addr_of_786_final_reg",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => array_obj_ref_785_root_address,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => arrayidx176_787,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1024_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1024_inst_req_0;
      type_cast_1024_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1024_inst_req_1;
      type_cast_1024_inst_ack_1<= rack(0);
      type_cast_1024_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1024_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp235x_xop_1021,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => iNsTr_60_1025,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1047_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1047_inst_req_0;
      type_cast_1047_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1047_inst_req_1;
      type_cast_1047_inst_ack_1<= rack(0);
      type_cast_1047_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1047_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext_1066,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1047_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1083_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_1083_inst_req_0;
      type_cast_1083_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_1083_inst_req_1;
      type_cast_1083_inst_ack_1<= rack(0);
      type_cast_1083_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1083_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ret_val_x_x_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_134_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_134_inst_req_0;
      type_cast_134_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_134_inst_req_1;
      type_cast_134_inst_ack_1<= rack(0);
      type_cast_134_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_134_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3_131,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4_135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_146_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_146_inst_req_0;
      type_cast_146_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_146_inst_req_1;
      type_cast_146_inst_ack_1<= rack(0);
      type_cast_146_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_146_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_146_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_153_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_153_inst_req_0;
      type_cast_153_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_153_inst_req_1;
      type_cast_153_inst_ack_1<= rack(0);
      type_cast_153_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_153_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_153_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_155_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_155_inst_req_0;
      type_cast_155_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_155_inst_req_1;
      type_cast_155_inst_ack_1<= rack(0);
      type_cast_155_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_155_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4x_xlcssa1_143,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_155_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_185_inst_req_0;
      type_cast_185_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_185_inst_req_1;
      type_cast_185_inst_ack_1<= rack(0);
      type_cast_185_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp265_223,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_185_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_198_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_198_inst_req_0;
      type_cast_198_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_198_inst_req_1;
      type_cast_198_inst_ack_1<= rack(0);
      type_cast_198_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_198_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp3_195,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc22_199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_212_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_212_inst_req_0;
      type_cast_212_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_212_inst_req_1;
      type_cast_212_inst_ack_1<= rack(0);
      type_cast_212_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_212_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call15_209,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv16_213,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_253_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_253_inst_req_0;
      type_cast_253_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_253_inst_req_1;
      type_cast_253_inst_ack_1<= rack(0);
      type_cast_253_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_253_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29217_250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30218_254,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_263_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_263_inst_req_0;
      type_cast_263_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_263_inst_req_1;
      type_cast_263_inst_ack_1<= rack(0);
      type_cast_263_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_263_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext261_292,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_263_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_267_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_267_inst_req_0;
      type_cast_267_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_267_inst_req_1;
      type_cast_267_inst_ack_1<= rack(0);
      type_cast_267_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_267_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30218_254,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_267_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_269_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_269_inst_req_0;
      type_cast_269_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_269_inst_req_1;
      type_cast_269_inst_ack_1<= rack(0);
      type_cast_269_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_269_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_269_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_285_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_285_inst_req_0;
      type_cast_285_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_285_inst_req_1;
      type_cast_285_inst_ack_1<= rack(0);
      type_cast_285_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_285_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call29_282,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv30_286,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_309_inst_req_0;
      type_cast_309_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_309_inst_req_1;
      type_cast_309_inst_ack_1<= rack(0);
      type_cast_309_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 16,
        out_data_width => 16,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv30_286,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_309_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_319_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_319_inst_req_0;
      type_cast_319_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_319_inst_req_1;
      type_cast_319_inst_ack_1<= rack(0);
      type_cast_319_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_319_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call40_316,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv41_320,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_338_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_338_inst_req_0;
      type_cast_338_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_338_inst_req_1;
      type_cast_338_inst_ack_1<= rack(0);
      type_cast_338_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_338_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call42_335,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv43_339,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_357_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_357_inst_req_0;
      type_cast_357_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_357_inst_req_1;
      type_cast_357_inst_ack_1<= rack(0);
      type_cast_357_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_357_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call44_354,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv45_358,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_38_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_38_inst_req_0;
      type_cast_38_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_38_inst_req_1;
      type_cast_38_inst_ack_1<= rack(0);
      type_cast_38_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_38_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_35,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv_39,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_419_inst_req_0;
      type_cast_419_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_419_inst_req_1;
      type_cast_419_inst_ack_1<= rack(0);
      type_cast_419_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_419_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul50_416,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv51_420,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_486_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_486_inst_req_0;
      type_cast_486_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_486_inst_req_1;
      type_cast_486_inst_ack_1<= rack(0);
      type_cast_486_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_486_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => mul59_483,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv60_487,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_540_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_540_inst_req_0;
      type_cast_540_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_540_inst_req_1;
      type_cast_540_inst_ack_1<= rack(0);
      type_cast_540_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_540_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp6_537,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp7_541,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_569_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_569_inst_req_0;
      type_cast_569_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_569_inst_req_1;
      type_cast_569_inst_ack_1<= rack(0);
      type_cast_569_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_569_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext251_720,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_569_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_583_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_583_inst_req_0;
      type_cast_583_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_583_inst_req_1;
      type_cast_583_inst_ack_1<= rack(0);
      type_cast_583_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_583_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call69_580,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv70_584,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_596_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_596_inst_req_0;
      type_cast_596_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_596_inst_req_1;
      type_cast_596_inst_ack_1<= rack(0);
      type_cast_596_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_596_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call72_593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv74_597,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_614_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_614_inst_req_1;
      type_cast_614_inst_ack_1<= rack(0);
      type_cast_614_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_614_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call77_611,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv79_615,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_62_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_62_inst_req_0;
      type_cast_62_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_62_inst_req_1;
      type_cast_62_inst_ack_1<= rack(0);
      type_cast_62_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_62_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call3228_59,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv4229_63,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_632_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_632_inst_req_0;
      type_cast_632_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_632_inst_req_1;
      type_cast_632_inst_ack_1<= rack(0);
      type_cast_632_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_632_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call83_629,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv85_633,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_650_inst_req_0;
      type_cast_650_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_650_inst_req_1;
      type_cast_650_inst_ack_1<= rack(0);
      type_cast_650_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_650_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call89_647,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv91_651,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_668_inst_req_0;
      type_cast_668_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_668_inst_req_1;
      type_cast_668_inst_ack_1<= rack(0);
      type_cast_668_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_668_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call95_665,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv97_669,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_686_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_686_inst_req_0;
      type_cast_686_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_686_inst_req_1;
      type_cast_686_inst_ack_1<= rack(0);
      type_cast_686_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_686_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call101_683,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv103_687,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_704_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_704_inst_req_0;
      type_cast_704_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_704_inst_req_1;
      type_cast_704_inst_ack_1<= rack(0);
      type_cast_704_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_704_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call107_701,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv109_705,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_750_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_750_inst_req_0;
      type_cast_750_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_750_inst_req_1;
      type_cast_750_inst_ack_1<= rack(0);
      type_cast_750_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_750_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp14_747,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tmp15_751,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_76_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_76_inst_req_0;
      type_cast_76_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_76_inst_req_1;
      type_cast_76_inst_ack_1<= rack(0);
      type_cast_76_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_76_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp270_113,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_76_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_779_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_779_inst_req_0;
      type_cast_779_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_779_inst_req_1;
      type_cast_779_inst_ack_1<= rack(0);
      type_cast_779_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_779_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => indvarx_xnext241_930,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_779_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_793_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_793_inst_req_0;
      type_cast_793_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_793_inst_req_1;
      type_cast_793_inst_ack_1<= rack(0);
      type_cast_793_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_793_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call129_790,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv130_794,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_806_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_806_inst_req_0;
      type_cast_806_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_806_inst_req_1;
      type_cast_806_inst_ack_1<= rack(0);
      type_cast_806_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_806_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call133_803,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv135_807,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_824_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_824_inst_req_0;
      type_cast_824_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_824_inst_req_1;
      type_cast_824_inst_ack_1<= rack(0);
      type_cast_824_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_824_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call139_821,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv141_825,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_83_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_83_inst_req_0;
      type_cast_83_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_83_inst_req_1;
      type_cast_83_inst_ack_1<= rack(0);
      type_cast_83_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_83_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4_135,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_83_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_842_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_842_inst_req_0;
      type_cast_842_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_842_inst_req_1;
      type_cast_842_inst_ack_1<= rack(0);
      type_cast_842_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_842_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call145_839,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv147_843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_85_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_85_inst_req_0;
      type_cast_85_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_85_inst_req_1;
      type_cast_85_inst_ack_1<= rack(0);
      type_cast_85_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_85_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => conv4229_63,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_85_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_860_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_860_inst_req_0;
      type_cast_860_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_860_inst_req_1;
      type_cast_860_inst_ack_1<= rack(0);
      type_cast_860_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_860_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call151_857,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv153_861,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_878_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_878_inst_req_0;
      type_cast_878_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_878_inst_req_1;
      type_cast_878_inst_ack_1<= rack(0);
      type_cast_878_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_878_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call157_875,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv159_879,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_896_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_896_inst_req_0;
      type_cast_896_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_896_inst_req_1;
      type_cast_896_inst_ack_1<= rack(0);
      type_cast_896_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_896_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call163_893,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv165_897,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_914_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_914_inst_req_0;
      type_cast_914_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_914_inst_req_1;
      type_cast_914_inst_ack_1<= rack(0);
      type_cast_914_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_914_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call169_911,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => conv171_915,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_95_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= type_cast_95_inst_req_0;
      type_cast_95_inst_ack_0<= wack(0);
      rreq(0) <= type_cast_95_inst_req_1;
      type_cast_95_inst_ack_1<= rack(0);
      type_cast_95_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_95_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tmp_92,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inc_96,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence STORE_padding_311_gather_scatter
    process(conv30x_xlcssa_306) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30x_xlcssa_306;
      ov(15 downto 0) := iv;
      STORE_padding_311_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_rename
    process(R_indvar268_100_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar268_100_resized;
      ov(6 downto 0) := iv;
      R_indvar268_100_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_index_1_resize
    process(indvar268_73) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar268_73;
      ov := iv(6 downto 0);
      R_indvar268_100_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_101_root_address_inst
    process(array_obj_ref_101_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_101_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_101_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1053_index_1_rename
    process(R_indvar_1052_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar_1052_resized;
      ov(13 downto 0) := iv;
      R_indvar_1052_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1053_index_1_resize
    process(indvar_1041) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar_1041;
      ov := iv(13 downto 0);
      R_indvar_1052_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1053_root_address_inst
    process(array_obj_ref_1053_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1053_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_1053_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_index_1_rename
    process(R_indvar263_203_resized) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar263_203_resized;
      ov(6 downto 0) := iv;
      R_indvar263_203_scaled <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_index_1_resize
    process(indvar263_182) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar263_182;
      ov := iv(6 downto 0);
      R_indvar263_203_resized <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_204_root_address_inst
    process(array_obj_ref_204_final_offset) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_204_final_offset;
      ov(6 downto 0) := iv;
      array_obj_ref_204_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_0_rename
    process(R_indvar260_272_resized) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_272_resized;
      ov(0 downto 0) := iv;
      R_indvar260_272_scaled <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_0_resize
    process(indvar260_257) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar260_257;
      ov := iv(0 downto 0);
      R_indvar260_272_resized <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_index_offset
    process(R_indvar260_272_scaled) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar260_272_scaled;
      ov(0 downto 0) := iv;
      array_obj_ref_273_final_offset <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_273_root_address_inst
    process(array_obj_ref_273_final_offset) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_273_final_offset;
      ov(0 downto 0) := iv;
      array_obj_ref_273_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_index_1_rename
    process(R_indvar250_574_resized) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar250_574_resized;
      ov(13 downto 0) := iv;
      R_indvar250_574_scaled <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_index_1_resize
    process(indvar250_563) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar250_563;
      ov := iv(13 downto 0);
      R_indvar250_574_resized <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_575_root_address_inst
    process(array_obj_ref_575_final_offset) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_575_final_offset;
      ov(13 downto 0) := iv;
      array_obj_ref_575_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_index_1_rename
    process(R_indvar240_784_resized) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_indvar240_784_resized;
      ov(10 downto 0) := iv;
      R_indvar240_784_scaled <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_index_1_resize
    process(indvar240_773) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := indvar240_773;
      ov := iv(10 downto 0);
      R_indvar240_784_resized <= ov(10 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_785_root_address_inst
    process(array_obj_ref_785_final_offset) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_785_final_offset;
      ov(10 downto 0) := iv;
      array_obj_ref_785_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1057_addr_0
    process(ptr_deref_1057_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1057_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_1057_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1057_base_resize
    process(arrayidx196_1055) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx196_1055;
      ov := iv(13 downto 0);
      ptr_deref_1057_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1057_gather_scatter
    process(type_cast_1059_wire_constant) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_1059_wire_constant;
      ov(63 downto 0) := iv;
      ptr_deref_1057_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_1057_root_address_inst
    process(ptr_deref_1057_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_1057_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_1057_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_addr_0
    process(ptr_deref_105_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_base_resize
    process(arrayidx_103) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx_103;
      ov := iv(6 downto 0);
      ptr_deref_105_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_gather_scatter
    process(conv4231_80) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4231_80;
      ov(31 downto 0) := iv;
      ptr_deref_105_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_105_root_address_inst
    process(ptr_deref_105_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_105_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_105_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_addr_0
    process(ptr_deref_122_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_base_resize
    process(iNsTr_13_119) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_13_119;
      ov := iv(6 downto 0);
      ptr_deref_122_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_gather_scatter
    process(ptr_deref_122_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_data_0;
      ov(31 downto 0) := iv;
      tmp1_123 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_122_root_address_inst
    process(ptr_deref_122_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_122_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_122_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_addr_0
    process(ptr_deref_164_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_164_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_164_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_base_resize
    process(iNsTr_5_162) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_5_162;
      ov := iv(6 downto 0);
      ptr_deref_164_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_gather_scatter
    process(conv4x_xlcssa_150) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv4x_xlcssa_150;
      ov(31 downto 0) := iv;
      ptr_deref_164_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_164_root_address_inst
    process(ptr_deref_164_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_164_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_164_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_addr_0
    process(ptr_deref_215_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_215_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_215_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_base_resize
    process(arrayidx19_206) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx19_206;
      ov := iv(6 downto 0);
      ptr_deref_215_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_gather_scatter
    process(conv16_213) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv16_213;
      ov(31 downto 0) := iv;
      ptr_deref_215_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_215_root_address_inst
    process(ptr_deref_215_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_215_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_215_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_addr_0
    process(ptr_deref_232_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_232_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_base_resize
    process(iNsTr_21_229) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_21_229;
      ov := iv(6 downto 0);
      ptr_deref_232_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_gather_scatter
    process(ptr_deref_232_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_data_0;
      ov(31 downto 0) := iv;
      tmp11_233 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_232_root_address_inst
    process(ptr_deref_232_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_232_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_232_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_addr_0
    process(ptr_deref_277_root_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_277_root_address;
      ov(0 downto 0) := iv;
      ptr_deref_277_word_address_0 <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_base_resize
    process(arrayidx33_275) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx33_275;
      ov := iv(0 downto 0);
      ptr_deref_277_resized_base_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_gather_scatter
    process(conv30220_264) --
      variable iv : std_logic_vector(15 downto 0);
      variable ov : std_logic_vector(15 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv30220_264;
      ov(15 downto 0) := iv;
      ptr_deref_277_data_0 <= ov(15 downto 0);
      --
    end process;
    -- equivalence ptr_deref_277_root_address_inst
    process(ptr_deref_277_resized_base_address) --
      variable iv : std_logic_vector(0 downto 0);
      variable ov : std_logic_vector(0 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_277_resized_base_address;
      ov(0 downto 0) := iv;
      ptr_deref_277_root_address <= ov(0 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_addr_0
    process(ptr_deref_330_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_330_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_330_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_base_resize
    process(iNsTr_26_328) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_26_328;
      ov := iv(6 downto 0);
      ptr_deref_330_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_gather_scatter
    process(conv41_320) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv41_320;
      ov(31 downto 0) := iv;
      ptr_deref_330_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_330_root_address_inst
    process(ptr_deref_330_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_330_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_330_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_addr_0
    process(ptr_deref_349_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_349_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_base_resize
    process(iNsTr_29_347) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_29_347;
      ov := iv(6 downto 0);
      ptr_deref_349_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_gather_scatter
    process(conv43_339) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv43_339;
      ov(31 downto 0) := iv;
      ptr_deref_349_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_349_root_address_inst
    process(ptr_deref_349_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_349_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_349_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_addr_0
    process(ptr_deref_368_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_368_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_368_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_base_resize
    process(iNsTr_32_366) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_32_366;
      ov := iv(6 downto 0);
      ptr_deref_368_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_gather_scatter
    process(conv45_358) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv45_358;
      ov(31 downto 0) := iv;
      ptr_deref_368_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_368_root_address_inst
    process(ptr_deref_368_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_368_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_368_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_addr_0
    process(ptr_deref_381_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_base_resize
    process(iNsTr_34_378) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_34_378;
      ov := iv(6 downto 0);
      ptr_deref_381_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_gather_scatter
    process(ptr_deref_381_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_data_0;
      ov(31 downto 0) := iv;
      tmp47_382 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_381_root_address_inst
    process(ptr_deref_381_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_381_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_381_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_addr_0
    process(ptr_deref_393_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_393_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_base_resize
    process(iNsTr_35_390) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_35_390;
      ov := iv(6 downto 0);
      ptr_deref_393_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_gather_scatter
    process(ptr_deref_393_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_data_0;
      ov(31 downto 0) := iv;
      tmp48_394 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_393_root_address_inst
    process(ptr_deref_393_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_393_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_393_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_addr_0
    process(ptr_deref_405_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_405_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_base_resize
    process(iNsTr_36_402) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_36_402;
      ov := iv(6 downto 0);
      ptr_deref_405_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_gather_scatter
    process(ptr_deref_405_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_data_0;
      ov(31 downto 0) := iv;
      tmp49_406 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_405_root_address_inst
    process(ptr_deref_405_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_405_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_405_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_addr_0
    process(ptr_deref_431_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_431_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_base_resize
    process(iNsTr_37_428) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_37_428;
      ov := iv(6 downto 0);
      ptr_deref_431_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_gather_scatter
    process(ptr_deref_431_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_data_0;
      ov(31 downto 0) := iv;
      tmp53_432 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_431_root_address_inst
    process(ptr_deref_431_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_431_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_431_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_addr_0
    process(ptr_deref_443_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_443_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_base_resize
    process(iNsTr_38_440) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_38_440;
      ov := iv(6 downto 0);
      ptr_deref_443_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_gather_scatter
    process(ptr_deref_443_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_data_0;
      ov(31 downto 0) := iv;
      tmp54_444 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_443_root_address_inst
    process(ptr_deref_443_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_443_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_443_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_addr_0
    process(ptr_deref_455_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_455_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_base_resize
    process(iNsTr_39_452) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_39_452;
      ov := iv(6 downto 0);
      ptr_deref_455_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_gather_scatter
    process(ptr_deref_455_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_data_0;
      ov(31 downto 0) := iv;
      tmp56_456 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_455_root_address_inst
    process(ptr_deref_455_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_455_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_455_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_addr_0
    process(ptr_deref_467_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_467_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_base_resize
    process(iNsTr_40_464) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_40_464;
      ov := iv(6 downto 0);
      ptr_deref_467_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_gather_scatter
    process(ptr_deref_467_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_data_0;
      ov(31 downto 0) := iv;
      tmp58_468 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_467_root_address_inst
    process(ptr_deref_467_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_467_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_467_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_addr_0
    process(ptr_deref_47_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_base_resize
    process(iNsTr_1_45) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_1_45;
      ov := iv(6 downto 0);
      ptr_deref_47_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_gather_scatter
    process(conv_39) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := conv_39;
      ov(31 downto 0) := iv;
      ptr_deref_47_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_47_root_address_inst
    process(ptr_deref_47_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_47_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_47_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_addr_0
    process(ptr_deref_712_root_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_712_root_address;
      ov(13 downto 0) := iv;
      ptr_deref_712_word_address_0 <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_base_resize
    process(arrayidx114_577) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx114_577;
      ov := iv(13 downto 0);
      ptr_deref_712_resized_base_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_gather_scatter
    process(add110_710) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add110_710;
      ov(63 downto 0) := iv;
      ptr_deref_712_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_712_root_address_inst
    process(ptr_deref_712_resized_base_address) --
      variable iv : std_logic_vector(13 downto 0);
      variable ov : std_logic_vector(13 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_712_resized_base_address;
      ov(13 downto 0) := iv;
      ptr_deref_712_root_address <= ov(13 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_addr_0
    process(ptr_deref_922_root_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_922_root_address;
      ov(10 downto 0) := iv;
      ptr_deref_922_word_address_0 <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_base_resize
    process(arrayidx176_787) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := arrayidx176_787;
      ov := iv(10 downto 0);
      ptr_deref_922_resized_base_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_gather_scatter
    process(add172_920) --
      variable iv : std_logic_vector(63 downto 0);
      variable ov : std_logic_vector(63 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := add172_920;
      ov(63 downto 0) := iv;
      ptr_deref_922_data_0 <= ov(63 downto 0);
      --
    end process;
    -- equivalence ptr_deref_922_root_address_inst
    process(ptr_deref_922_resized_base_address) --
      variable iv : std_logic_vector(10 downto 0);
      variable ov : std_logic_vector(10 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_922_resized_base_address;
      ov(10 downto 0) := iv;
      ptr_deref_922_root_address <= ov(10 downto 0);
      --
    end process;
    -- equivalence ptr_deref_955_addr_0
    process(ptr_deref_955_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_955_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_955_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_955_base_resize
    process(iNsTr_45_952) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_45_952;
      ov := iv(6 downto 0);
      ptr_deref_955_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_955_gather_scatter
    process(ptr_deref_955_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_955_data_0;
      ov(31 downto 0) := iv;
      tmp182_956 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_955_root_address_inst
    process(ptr_deref_955_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_955_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_955_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_967_addr_0
    process(ptr_deref_967_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_967_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_967_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_967_base_resize
    process(iNsTr_46_964) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_46_964;
      ov := iv(6 downto 0);
      ptr_deref_967_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_967_gather_scatter
    process(ptr_deref_967_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_967_data_0;
      ov(31 downto 0) := iv;
      tmp183_968 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_967_root_address_inst
    process(ptr_deref_967_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_967_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_967_root_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_979_addr_0
    process(ptr_deref_979_root_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_979_root_address;
      ov(6 downto 0) := iv;
      ptr_deref_979_word_address_0 <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_979_base_resize
    process(iNsTr_47_976) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := iNsTr_47_976;
      ov := iv(6 downto 0);
      ptr_deref_979_resized_base_address <= ov(6 downto 0);
      --
    end process;
    -- equivalence ptr_deref_979_gather_scatter
    process(ptr_deref_979_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_979_data_0;
      ov(31 downto 0) := iv;
      tmp185_980 <= ov(31 downto 0);
      --
    end process;
    -- equivalence ptr_deref_979_root_address_inst
    process(ptr_deref_979_resized_base_address) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(6 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := ptr_deref_979_resized_base_address;
      ov(6 downto 0) := iv;
      ptr_deref_979_root_address <= ov(6 downto 0);
      --
    end process;
    if_stmt_1072_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond20_1071;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1072_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1072_branch_req_0,
          ack0 => if_stmt_1072_branch_ack_0,
          ack1 => if_stmt_1072_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_136_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp_128;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_136_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_136_branch_req_0,
          ack0 => if_stmt_136_branch_ack_0,
          ack1 => if_stmt_136_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_173_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12223_172;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_173_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_173_branch_req_0,
          ack0 => if_stmt_173_branch_ack_0,
          ack1 => if_stmt_173_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_239_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp12_238;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_239_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_239_branch_req_0,
          ack0 => if_stmt_239_branch_ack_0,
          ack1 => if_stmt_239_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_299_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_298;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_299_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_299_branch_req_0,
          ack0 => if_stmt_299_branch_ack_0,
          ack1 => if_stmt_299_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_500_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp65213_499;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_500_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_500_branch_req_0,
          ack0 => if_stmt_500_branch_ack_0,
          ack1 => if_stmt_500_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_521_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp124208_520;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_521_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_521_branch_req_0,
          ack0 => if_stmt_521_branch_ack_0,
          ack1 => if_stmt_521_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_64_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp227_56;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_64_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_64_branch_req_0,
          ack0 => if_stmt_64_branch_ack_0,
          ack1 => if_stmt_64_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_726_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond10_725;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_726_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_726_branch_req_0,
          ack0 => if_stmt_726_branch_ack_0,
          ack1 => if_stmt_726_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_936_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond19_935;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_936_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_936_branch_req_0,
          ack0 => if_stmt_936_branch_ack_0,
          ack1 => if_stmt_936_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_997_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= cmp191204_996;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_997_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_997_branch_req_0,
          ack0 => if_stmt_997_branch_ack_0,
          ack1 => if_stmt_997_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_1020_inst
    process(tmp235_1009) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(tmp235_1009, type_cast_1019_wire_constant, tmp_var);
      tmp235x_xop_1021 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1030_inst
    process(iNsTr_60_1025) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(iNsTr_60_1025, type_cast_1029_wire_constant, tmp_var);
      xx_xop_1031 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_1065_inst
    process(indvar_1041) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar_1041, type_cast_1064_wire_constant, tmp_var);
      indvarx_xnext_1066 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_112_inst
    process(indvar268_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_73, type_cast_111_wire_constant, tmp_var);
      tmp270_113 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_194_inst
    process(indvar263_182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_182, type_cast_193_wire_constant, tmp_var);
      tmp3_195 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_222_inst
    process(indvar263_182) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar263_182, type_cast_221_wire_constant, tmp_var);
      tmp265_223 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_291_inst
    process(indvar260_257) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar260_257, type_cast_290_wire_constant, tmp_var);
      indvarx_xnext261_292 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_719_inst
    process(indvar250_563) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar250_563, type_cast_718_wire_constant, tmp_var);
      indvarx_xnext251_720 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_91_inst
    process(indvar268_73) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar268_73, type_cast_90_wire_constant, tmp_var);
      tmp_92 <= tmp_var; --
    end process;
    -- binary operator ADD_u64_u64_929_inst
    process(indvar240_773) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAdd_proc(indvar240_773, type_cast_928_wire_constant, tmp_var);
      indvarx_xnext241_930 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_492_inst
    process(conv51_420) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv51_420, type_cast_491_wire_constant, tmp_var);
      shr212x_xmask_493 <= tmp_var; --
    end process;
    -- binary operator AND_u64_u64_513_inst
    process(conv60_487) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntAnd_proc(conv60_487, type_cast_512_wire_constant, tmp_var);
      shr123207x_xmask_514 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_171_inst
    process(conv4x_xlcssa_150) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(conv4x_xlcssa_150, type_cast_170_wire_constant, tmp_var);
      cmp12223_172 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1070_inst
    process(indvarx_xnext_1066, tmp239_1038) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext_1066, tmp239_1038, tmp_var);
      exitcond20_1071 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_297_inst
    process(indvarx_xnext261_292) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext261_292, type_cast_296_wire_constant, tmp_var);
      exitcond_298 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_498_inst
    process(shr212x_xmask_493) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr212x_xmask_493, type_cast_497_wire_constant, tmp_var);
      cmp65213_499 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_519_inst
    process(shr123207x_xmask_514) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shr123207x_xmask_514, type_cast_518_wire_constant, tmp_var);
      cmp124208_520 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_724_inst
    process(indvarx_xnext251_720, umax_560) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext251_720, umax_560, tmp_var);
      exitcond10_725 <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_934_inst
    process(indvarx_xnext241_930, umax18_770) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(indvarx_xnext241_930, umax18_770, tmp_var);
      exitcond19_935 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_54_inst
    process(call_35) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(call_35, type_cast_53_wire_constant, tmp_var);
      cmp227_56 <= tmp_var; --
    end process;
    -- binary operator LSHR_u32_u32_1008_inst
    process(mul186_990) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(mul186_990, type_cast_1007_wire_constant, tmp_var);
      tmp235_1009 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_546_inst
    process(tmp7_541) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp7_541, type_cast_545_wire_constant, tmp_var);
      tmp8_547 <= tmp_var; --
    end process;
    -- binary operator LSHR_u64_u64_756_inst
    process(tmp15_751) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntLSHR_proc(tmp15_751, type_cast_755_wire_constant, tmp_var);
      tmp16_757 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_410_inst
    process(tmp48_394, tmp47_382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_394, tmp47_382, tmp_var);
      mul_411 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_415_inst
    process(mul_411, tmp49_406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul_411, tmp49_406, tmp_var);
      mul50_416 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_472_inst
    process(tmp54_444, tmp53_432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_444, tmp53_432, tmp_var);
      mul55_473 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_477_inst
    process(mul55_473, tmp56_456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul55_473, tmp56_456, tmp_var);
      mul57_478 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_482_inst
    process(mul57_478, tmp58_468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul57_478, tmp58_468, tmp_var);
      mul59_483 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_531_inst
    process(tmp48_394, tmp47_382) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp48_394, tmp47_382, tmp_var);
      tmp5_532 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_536_inst
    process(tmp5_532, tmp49_406) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp5_532, tmp49_406, tmp_var);
      tmp6_537 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_736_inst
    process(tmp54_444, tmp53_432) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp54_444, tmp53_432, tmp_var);
      tmp12_737 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_741_inst
    process(tmp12_737, tmp56_456) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp12_737, tmp56_456, tmp_var);
      tmp13_742 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_746_inst
    process(tmp13_742, tmp58_468) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp13_742, tmp58_468, tmp_var);
      tmp14_747 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_984_inst
    process(tmp183_968, tmp182_956) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(tmp183_968, tmp182_956, tmp_var);
      mul184_985 <= tmp_var; --
    end process;
    -- binary operator MUL_u32_u32_989_inst
    process(mul184_985, tmp185_980) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntMul_proc(mul184_985, tmp185_980, tmp_var);
      mul186_990 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_601_inst
    process(shl_590, conv74_597) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl_590, conv74_597, tmp_var);
      add_602 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_619_inst
    process(shl76_608, conv79_615) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl76_608, conv79_615, tmp_var);
      add80_620 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_637_inst
    process(shl82_626, conv85_633) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl82_626, conv85_633, tmp_var);
      add86_638 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_655_inst
    process(shl88_644, conv91_651) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl88_644, conv91_651, tmp_var);
      add92_656 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_673_inst
    process(shl94_662, conv97_669) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl94_662, conv97_669, tmp_var);
      add98_674 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_691_inst
    process(shl100_680, conv103_687) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl100_680, conv103_687, tmp_var);
      add104_692 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_709_inst
    process(shl106_698, conv109_705) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl106_698, conv109_705, tmp_var);
      add110_710 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_811_inst
    process(shl132_800, conv135_807) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl132_800, conv135_807, tmp_var);
      add136_812 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_829_inst
    process(shl138_818, conv141_825) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl138_818, conv141_825, tmp_var);
      add142_830 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_847_inst
    process(shl144_836, conv147_843) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl144_836, conv147_843, tmp_var);
      add148_848 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_865_inst
    process(shl150_854, conv153_861) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl150_854, conv153_861, tmp_var);
      add154_866 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_883_inst
    process(shl156_872, conv159_879) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl156_872, conv159_879, tmp_var);
      add160_884 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_901_inst
    process(shl162_890, conv165_897) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl162_890, conv165_897, tmp_var);
      add166_902 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_919_inst
    process(shl168_908, conv171_915) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(shl168_908, conv171_915, tmp_var);
      add172_920 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_589_inst
    process(conv70_584) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv70_584, type_cast_588_wire_constant, tmp_var);
      shl_590 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_607_inst
    process(add_602) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add_602, type_cast_606_wire_constant, tmp_var);
      shl76_608 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_625_inst
    process(add80_620) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add80_620, type_cast_624_wire_constant, tmp_var);
      shl82_626 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_643_inst
    process(add86_638) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add86_638, type_cast_642_wire_constant, tmp_var);
      shl88_644 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_661_inst
    process(add92_656) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add92_656, type_cast_660_wire_constant, tmp_var);
      shl94_662 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_679_inst
    process(add98_674) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add98_674, type_cast_678_wire_constant, tmp_var);
      shl100_680 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_697_inst
    process(add104_692) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add104_692, type_cast_696_wire_constant, tmp_var);
      shl106_698 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_799_inst
    process(conv130_794) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(conv130_794, type_cast_798_wire_constant, tmp_var);
      shl132_800 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_817_inst
    process(add136_812) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add136_812, type_cast_816_wire_constant, tmp_var);
      shl138_818 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_835_inst
    process(add142_830) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add142_830, type_cast_834_wire_constant, tmp_var);
      shl144_836 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_853_inst
    process(add148_848) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add148_848, type_cast_852_wire_constant, tmp_var);
      shl150_854 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_871_inst
    process(add154_866) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add154_866, type_cast_870_wire_constant, tmp_var);
      shl156_872 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_889_inst
    process(add160_884) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add160_884, type_cast_888_wire_constant, tmp_var);
      shl162_890 <= tmp_var; --
    end process;
    -- binary operator SHL_u64_u64_907_inst
    process(add166_902) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntSHL_proc(add166_902, type_cast_906_wire_constant, tmp_var);
      shl168_908 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1014_inst
    process(tmp235_1009) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp235_1009, type_cast_1013_wire_constant, tmp_var);
      tmp236_1015 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_995_inst
    process(mul186_990) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(mul186_990, type_cast_994_wire_constant, tmp_var);
      cmp191204_996 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_552_inst
    process(tmp8_547) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp8_547, type_cast_551_wire_constant, tmp_var);
      tmp9_553 <= tmp_var; --
    end process;
    -- binary operator UGT_u64_u1_762_inst
    process(tmp16_757) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tmp16_757, type_cast_761_wire_constant, tmp_var);
      tmp17_763 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_127_inst
    process(inc_96, tmp1_123) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc_96, tmp1_123, tmp_var);
      cmp_128 <= tmp_var; --
    end process;
    -- binary operator ULT_u32_u1_237_inst
    process(inc22_199, tmp11_233) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(inc22_199, tmp11_233, tmp_var);
      cmp12_238 <= tmp_var; --
    end process;
    -- shared split operator group (69) : array_obj_ref_101_index_offset 
    ApIntAdd_group_69: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar268_100_scaled;
      array_obj_ref_101_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_101_index_offset_req_0;
      array_obj_ref_101_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_101_index_offset_req_1;
      array_obj_ref_101_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_69_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_69_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_69",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : array_obj_ref_1053_index_offset 
    ApIntAdd_group_70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar_1052_scaled;
      array_obj_ref_1053_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_1053_index_offset_req_0;
      array_obj_ref_1053_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_1053_index_offset_req_1;
      array_obj_ref_1053_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_70_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_70_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_70",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : array_obj_ref_204_index_offset 
    ApIntAdd_group_71: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(6 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar263_203_scaled;
      array_obj_ref_204_final_offset <= data_out(6 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_204_index_offset_req_0;
      array_obj_ref_204_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_204_index_offset_req_1;
      array_obj_ref_204_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_71_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_71_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_71",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 7,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 7,
          constant_operand => "0000010",
          constant_width => 7,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : array_obj_ref_575_index_offset 
    ApIntAdd_group_72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar250_574_scaled;
      array_obj_ref_575_final_offset <= data_out(13 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_575_index_offset_req_0;
      array_obj_ref_575_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_575_index_offset_req_1;
      array_obj_ref_575_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_72_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_72_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_72",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : array_obj_ref_785_index_offset 
    ApIntAdd_group_73: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= R_indvar240_784_scaled;
      array_obj_ref_785_final_offset <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= array_obj_ref_785_index_offset_req_0;
      array_obj_ref_785_index_offset_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_785_index_offset_req_1;
      array_obj_ref_785_index_offset_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_73_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_73_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_73",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000100001",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared load operator group (0) : ptr_deref_122_load_0 ptr_deref_381_load_0 ptr_deref_393_load_0 ptr_deref_405_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= ptr_deref_122_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_381_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_393_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_405_load_0_req_0;
      ptr_deref_122_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_381_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_393_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_405_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_122_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_381_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_393_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_405_load_0_req_1;
      ptr_deref_122_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_381_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_393_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_405_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_122_word_address_0 & ptr_deref_381_word_address_0 & ptr_deref_393_word_address_0 & ptr_deref_405_word_address_0;
      ptr_deref_122_data_0 <= data_out(127 downto 96);
      ptr_deref_381_data_0 <= data_out(95 downto 64);
      ptr_deref_393_data_0 <= data_out(63 downto 32);
      ptr_deref_405_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 7,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_467_load_0 ptr_deref_431_load_0 ptr_deref_443_load_0 ptr_deref_455_load_0 ptr_deref_232_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(34 downto 0);
      signal data_out: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 4 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 4 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 4 downto 0);
      signal guard_vector : std_logic_vector( 4 downto 0);
      constant inBUFs : IntegerArray(4 downto 0) := (4 => 0, 3 => 0, 2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(4 downto 0) := (4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(4 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false);
      constant guardBuffering: IntegerArray(4 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2);
      -- 
    begin -- 
      reqL_unguarded(4) <= ptr_deref_467_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_431_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_443_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_455_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_232_load_0_req_0;
      ptr_deref_467_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_431_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_443_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_455_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_232_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(4) <= ptr_deref_467_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_431_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_443_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_455_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_232_load_0_req_1;
      ptr_deref_467_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_431_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_443_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_455_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_232_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      LoadGroup1_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup1_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup1_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup1_gI: SplitGuardInterface generic map(name => "LoadGroup1_gI", nreqs => 5, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_467_word_address_0 & ptr_deref_431_word_address_0 & ptr_deref_443_word_address_0 & ptr_deref_455_word_address_0 & ptr_deref_232_word_address_0;
      ptr_deref_467_data_0 <= data_out(159 downto 128);
      ptr_deref_431_data_0 <= data_out(127 downto 96);
      ptr_deref_443_data_0 <= data_out(95 downto 64);
      ptr_deref_455_data_0 <= data_out(63 downto 32);
      ptr_deref_232_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup1", addr_width => 7,
        num_reqs => 5,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup1 load-complete ",
        data_width => 32,
        num_reqs => 5,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_979_load_0 ptr_deref_967_load_0 ptr_deref_955_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(20 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_979_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_967_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_955_load_0_req_0;
      ptr_deref_979_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_967_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_955_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_979_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_967_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_955_load_0_req_1;
      ptr_deref_979_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_967_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_955_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      LoadGroup2_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup2_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup2_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup2_gI: SplitGuardInterface generic map(name => "LoadGroup2_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= ptr_deref_979_word_address_0 & ptr_deref_967_word_address_0 & ptr_deref_955_word_address_0;
      ptr_deref_979_data_0 <= data_out(95 downto 64);
      ptr_deref_967_data_0 <= data_out(63 downto 32);
      ptr_deref_955_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup2", addr_width => 7,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup2 load-complete ",
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared store operator group (0) : STORE_padding_311_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= STORE_padding_311_store_0_req_0;
      STORE_padding_311_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= STORE_padding_311_store_0_req_1;
      STORE_padding_311_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= STORE_padding_311_word_address_0;
      data_in <= STORE_padding_311_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(15 downto 0),
          mtag => memory_space_6_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1057_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_1057_store_0_req_0;
      ptr_deref_1057_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1057_store_0_req_1;
      ptr_deref_1057_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup1_gI: SplitGuardInterface generic map(name => "StoreGroup1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1057_word_address_0;
      data_in <= ptr_deref_1057_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup1 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(13 downto 0),
          mdata => memory_space_5_sr_data(63 downto 0),
          mtag => memory_space_5_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup1 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_47_store_0 ptr_deref_105_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_47_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_105_store_0_req_0;
      ptr_deref_47_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_105_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_47_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_105_store_0_req_1;
      ptr_deref_47_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_105_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup2_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup2_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup2_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup2_gI: SplitGuardInterface generic map(name => "StoreGroup2_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_47_word_address_0 & ptr_deref_105_word_address_0;
      data_in <= ptr_deref_47_data_0 & ptr_deref_105_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup2 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup2 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_164_store_0 ptr_deref_215_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_164_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_215_store_0_req_0;
      ptr_deref_164_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_215_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_164_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_215_store_0_req_1;
      ptr_deref_164_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_215_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      StoreGroup3_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup3_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup3_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup3_gI: SplitGuardInterface generic map(name => "StoreGroup3_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_164_word_address_0 & ptr_deref_215_word_address_0;
      data_in <= ptr_deref_164_data_0 & ptr_deref_215_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup3 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup3 Complete ",
          num_reqs => 2,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_277_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_277_store_0_req_0;
      ptr_deref_277_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_277_store_0_req_1;
      ptr_deref_277_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup4_gI: SplitGuardInterface generic map(name => "StoreGroup4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_277_word_address_0;
      data_in <= ptr_deref_277_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup4 Req ", addr_width => 1,
        data_width => 16,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(15 downto 0),
          mtag => memory_space_7_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup4 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_330_store_0 ptr_deref_349_store_0 ptr_deref_368_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(20 downto 0);
      signal data_in: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      constant inBUFs : IntegerArray(2 downto 0) := (2 => 0, 1 => 0, 0 => 0);
      constant outBUFs : IntegerArray(2 downto 0) := (2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(2 downto 0) := (0 => false, 1 => false, 2 => false);
      constant guardBuffering: IntegerArray(2 downto 0)  := (0 => 2, 1 => 2, 2 => 2);
      -- 
    begin -- 
      reqL_unguarded(2) <= ptr_deref_330_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_349_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_368_store_0_req_0;
      ptr_deref_330_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_349_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_368_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_330_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_349_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_368_store_0_req_1;
      ptr_deref_330_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_349_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_368_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      StoreGroup5_accessRegulator_0: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_1: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      StoreGroup5_accessRegulator_2: access_regulator_base generic map (name => "StoreGroup5_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      StoreGroup5_gI: SplitGuardInterface generic map(name => "StoreGroup5_gI", nreqs => 3, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_330_word_address_0 & ptr_deref_349_word_address_0 & ptr_deref_368_word_address_0;
      data_in <= ptr_deref_330_data_0 & ptr_deref_349_data_0 & ptr_deref_368_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup5 Req ", addr_width => 7,
        data_width => 32,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(19 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup5 Complete ",
          num_reqs => 3,
          detailed_buffering_per_output => outBUFs,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_712_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(13 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_712_store_0_req_0;
      ptr_deref_712_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_712_store_0_req_1;
      ptr_deref_712_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup6_gI: SplitGuardInterface generic map(name => "StoreGroup6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_712_word_address_0;
      data_in <= ptr_deref_712_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup6 Req ", addr_width => 14,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(63 downto 0),
          mtag => memory_space_3_sr_tag(18 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup6 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_922_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(10 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_922_store_0_req_0;
      ptr_deref_922_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_922_store_0_req_1;
      ptr_deref_922_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup7_gI: SplitGuardInterface generic map(name => "StoreGroup7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_922_word_address_0;
      data_in <= ptr_deref_922_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup7 Req ", addr_width => 11,
        data_width => 64,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 0,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(10 downto 0),
          mdata => memory_space_4_sr_data(63 downto 0),
          mtag => memory_space_4_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup7 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared inport operator group (0) : RPIPE_ConvTranspose_input_pipe_874_inst RPIPE_ConvTranspose_input_pipe_892_inst RPIPE_ConvTranspose_input_pipe_664_inst RPIPE_ConvTranspose_input_pipe_820_inst RPIPE_ConvTranspose_input_pipe_682_inst RPIPE_ConvTranspose_input_pipe_838_inst RPIPE_ConvTranspose_input_pipe_910_inst RPIPE_ConvTranspose_input_pipe_579_inst RPIPE_ConvTranspose_input_pipe_700_inst RPIPE_ConvTranspose_input_pipe_592_inst RPIPE_ConvTranspose_input_pipe_610_inst RPIPE_ConvTranspose_input_pipe_628_inst RPIPE_ConvTranspose_input_pipe_789_inst RPIPE_ConvTranspose_input_pipe_646_inst RPIPE_ConvTranspose_input_pipe_802_inst RPIPE_ConvTranspose_input_pipe_856_inst RPIPE_ConvTranspose_input_pipe_34_inst RPIPE_ConvTranspose_input_pipe_58_inst RPIPE_ConvTranspose_input_pipe_130_inst RPIPE_ConvTranspose_input_pipe_208_inst RPIPE_ConvTranspose_input_pipe_249_inst RPIPE_ConvTranspose_input_pipe_281_inst RPIPE_ConvTranspose_input_pipe_315_inst RPIPE_ConvTranspose_input_pipe_334_inst RPIPE_ConvTranspose_input_pipe_353_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(199 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 24 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 24 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 24 downto 0);
      signal guard_vector : std_logic_vector( 24 downto 0);
      constant outBUFs : IntegerArray(24 downto 0) := (24 => 1, 23 => 1, 22 => 1, 21 => 1, 20 => 1, 19 => 1, 18 => 1, 17 => 1, 16 => 1, 15 => 1, 14 => 1, 13 => 1, 12 => 1, 11 => 1, 10 => 1, 9 => 1, 8 => 1, 7 => 1, 6 => 1, 5 => 1, 4 => 1, 3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(24 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false, 4 => false, 5 => false, 6 => false, 7 => false, 8 => false, 9 => false, 10 => false, 11 => false, 12 => false, 13 => false, 14 => false, 15 => false, 16 => false, 17 => false, 18 => false, 19 => false, 20 => false, 21 => false, 22 => false, 23 => false, 24 => false);
      constant guardBuffering: IntegerArray(24 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2, 4 => 2, 5 => 2, 6 => 2, 7 => 2, 8 => 2, 9 => 2, 10 => 2, 11 => 2, 12 => 2, 13 => 2, 14 => 2, 15 => 2, 16 => 2, 17 => 2, 18 => 2, 19 => 2, 20 => 2, 21 => 2, 22 => 2, 23 => 2, 24 => 2);
      -- 
    begin -- 
      reqL_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_874_inst_req_0;
      reqL_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_892_inst_req_0;
      reqL_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_0;
      reqL_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_820_inst_req_0;
      reqL_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_0;
      reqL_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_838_inst_req_0;
      reqL_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_910_inst_req_0;
      reqL_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_0;
      reqL_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_0;
      reqL_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_592_inst_req_0;
      reqL_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_610_inst_req_0;
      reqL_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_628_inst_req_0;
      reqL_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_0;
      reqL_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_646_inst_req_0;
      reqL_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_802_inst_req_0;
      reqL_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_856_inst_req_0;
      reqL_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_0;
      reqL_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_0;
      reqL_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_130_inst_req_0;
      reqL_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_208_inst_req_0;
      reqL_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_249_inst_req_0;
      reqL_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_0;
      reqL_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_315_inst_req_0;
      reqL_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_334_inst_req_0;
      reqL_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_0;
      RPIPE_ConvTranspose_input_pipe_874_inst_ack_0 <= ackL_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_892_inst_ack_0 <= ackL_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_0 <= ackL_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_820_inst_ack_0 <= ackL_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_0 <= ackL_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_838_inst_ack_0 <= ackL_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_910_inst_ack_0 <= ackL_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_0 <= ackL_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_0 <= ackL_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_592_inst_ack_0 <= ackL_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_610_inst_ack_0 <= ackL_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_628_inst_ack_0 <= ackL_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_0 <= ackL_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_646_inst_ack_0 <= ackL_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_802_inst_ack_0 <= ackL_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_856_inst_ack_0 <= ackL_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_0 <= ackL_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_0 <= ackL_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_130_inst_ack_0 <= ackL_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_208_inst_ack_0 <= ackL_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_249_inst_ack_0 <= ackL_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_0 <= ackL_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_315_inst_ack_0 <= ackL_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_334_inst_ack_0 <= ackL_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(24) <= RPIPE_ConvTranspose_input_pipe_874_inst_req_1;
      reqR_unguarded(23) <= RPIPE_ConvTranspose_input_pipe_892_inst_req_1;
      reqR_unguarded(22) <= RPIPE_ConvTranspose_input_pipe_664_inst_req_1;
      reqR_unguarded(21) <= RPIPE_ConvTranspose_input_pipe_820_inst_req_1;
      reqR_unguarded(20) <= RPIPE_ConvTranspose_input_pipe_682_inst_req_1;
      reqR_unguarded(19) <= RPIPE_ConvTranspose_input_pipe_838_inst_req_1;
      reqR_unguarded(18) <= RPIPE_ConvTranspose_input_pipe_910_inst_req_1;
      reqR_unguarded(17) <= RPIPE_ConvTranspose_input_pipe_579_inst_req_1;
      reqR_unguarded(16) <= RPIPE_ConvTranspose_input_pipe_700_inst_req_1;
      reqR_unguarded(15) <= RPIPE_ConvTranspose_input_pipe_592_inst_req_1;
      reqR_unguarded(14) <= RPIPE_ConvTranspose_input_pipe_610_inst_req_1;
      reqR_unguarded(13) <= RPIPE_ConvTranspose_input_pipe_628_inst_req_1;
      reqR_unguarded(12) <= RPIPE_ConvTranspose_input_pipe_789_inst_req_1;
      reqR_unguarded(11) <= RPIPE_ConvTranspose_input_pipe_646_inst_req_1;
      reqR_unguarded(10) <= RPIPE_ConvTranspose_input_pipe_802_inst_req_1;
      reqR_unguarded(9) <= RPIPE_ConvTranspose_input_pipe_856_inst_req_1;
      reqR_unguarded(8) <= RPIPE_ConvTranspose_input_pipe_34_inst_req_1;
      reqR_unguarded(7) <= RPIPE_ConvTranspose_input_pipe_58_inst_req_1;
      reqR_unguarded(6) <= RPIPE_ConvTranspose_input_pipe_130_inst_req_1;
      reqR_unguarded(5) <= RPIPE_ConvTranspose_input_pipe_208_inst_req_1;
      reqR_unguarded(4) <= RPIPE_ConvTranspose_input_pipe_249_inst_req_1;
      reqR_unguarded(3) <= RPIPE_ConvTranspose_input_pipe_281_inst_req_1;
      reqR_unguarded(2) <= RPIPE_ConvTranspose_input_pipe_315_inst_req_1;
      reqR_unguarded(1) <= RPIPE_ConvTranspose_input_pipe_334_inst_req_1;
      reqR_unguarded(0) <= RPIPE_ConvTranspose_input_pipe_353_inst_req_1;
      RPIPE_ConvTranspose_input_pipe_874_inst_ack_1 <= ackR_unguarded(24);
      RPIPE_ConvTranspose_input_pipe_892_inst_ack_1 <= ackR_unguarded(23);
      RPIPE_ConvTranspose_input_pipe_664_inst_ack_1 <= ackR_unguarded(22);
      RPIPE_ConvTranspose_input_pipe_820_inst_ack_1 <= ackR_unguarded(21);
      RPIPE_ConvTranspose_input_pipe_682_inst_ack_1 <= ackR_unguarded(20);
      RPIPE_ConvTranspose_input_pipe_838_inst_ack_1 <= ackR_unguarded(19);
      RPIPE_ConvTranspose_input_pipe_910_inst_ack_1 <= ackR_unguarded(18);
      RPIPE_ConvTranspose_input_pipe_579_inst_ack_1 <= ackR_unguarded(17);
      RPIPE_ConvTranspose_input_pipe_700_inst_ack_1 <= ackR_unguarded(16);
      RPIPE_ConvTranspose_input_pipe_592_inst_ack_1 <= ackR_unguarded(15);
      RPIPE_ConvTranspose_input_pipe_610_inst_ack_1 <= ackR_unguarded(14);
      RPIPE_ConvTranspose_input_pipe_628_inst_ack_1 <= ackR_unguarded(13);
      RPIPE_ConvTranspose_input_pipe_789_inst_ack_1 <= ackR_unguarded(12);
      RPIPE_ConvTranspose_input_pipe_646_inst_ack_1 <= ackR_unguarded(11);
      RPIPE_ConvTranspose_input_pipe_802_inst_ack_1 <= ackR_unguarded(10);
      RPIPE_ConvTranspose_input_pipe_856_inst_ack_1 <= ackR_unguarded(9);
      RPIPE_ConvTranspose_input_pipe_34_inst_ack_1 <= ackR_unguarded(8);
      RPIPE_ConvTranspose_input_pipe_58_inst_ack_1 <= ackR_unguarded(7);
      RPIPE_ConvTranspose_input_pipe_130_inst_ack_1 <= ackR_unguarded(6);
      RPIPE_ConvTranspose_input_pipe_208_inst_ack_1 <= ackR_unguarded(5);
      RPIPE_ConvTranspose_input_pipe_249_inst_ack_1 <= ackR_unguarded(4);
      RPIPE_ConvTranspose_input_pipe_281_inst_ack_1 <= ackR_unguarded(3);
      RPIPE_ConvTranspose_input_pipe_315_inst_ack_1 <= ackR_unguarded(2);
      RPIPE_ConvTranspose_input_pipe_334_inst_ack_1 <= ackR_unguarded(1);
      RPIPE_ConvTranspose_input_pipe_353_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      guard_vector(12)  <=  '1';
      guard_vector(13)  <=  '1';
      guard_vector(14)  <=  '1';
      guard_vector(15)  <=  '1';
      guard_vector(16)  <=  '1';
      guard_vector(17)  <=  '1';
      guard_vector(18)  <=  '1';
      guard_vector(19)  <=  '1';
      guard_vector(20)  <=  '1';
      guard_vector(21)  <=  '1';
      guard_vector(22)  <=  '1';
      guard_vector(23)  <=  '1';
      guard_vector(24)  <=  '1';
      call157_875 <= data_out(199 downto 192);
      call163_893 <= data_out(191 downto 184);
      call95_665 <= data_out(183 downto 176);
      call139_821 <= data_out(175 downto 168);
      call101_683 <= data_out(167 downto 160);
      call145_839 <= data_out(159 downto 152);
      call169_911 <= data_out(151 downto 144);
      call69_580 <= data_out(143 downto 136);
      call107_701 <= data_out(135 downto 128);
      call72_593 <= data_out(127 downto 120);
      call77_611 <= data_out(119 downto 112);
      call83_629 <= data_out(111 downto 104);
      call129_790 <= data_out(103 downto 96);
      call89_647 <= data_out(95 downto 88);
      call133_803 <= data_out(87 downto 80);
      call151_857 <= data_out(79 downto 72);
      call_35 <= data_out(71 downto 64);
      call3228_59 <= data_out(63 downto 56);
      call3_131 <= data_out(55 downto 48);
      call15_209 <= data_out(47 downto 40);
      call29217_250 <= data_out(39 downto 32);
      call29_282 <= data_out(31 downto 24);
      call40_316 <= data_out(23 downto 16);
      call42_335 <= data_out(15 downto 8);
      call44_354 <= data_out(7 downto 0);
      ConvTranspose_input_pipe_read_0_gI: SplitGuardInterface generic map(name => "ConvTranspose_input_pipe_read_0_gI", nreqs => 25, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      ConvTranspose_input_pipe_read_0: InputPortRevised -- 
        generic map ( name => "ConvTranspose_input_pipe_read_0", data_width => 8,  num_reqs => 25,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => ConvTranspose_input_pipe_pipe_read_req(0),
          oack => ConvTranspose_input_pipe_pipe_read_ack(0),
          odata => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  -- 
end testConfigure_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    ConvTranspose_input_pipe_pipe_write_data: in std_logic_vector(7 downto 0);
    ConvTranspose_input_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    ConvTranspose_input_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_data: out std_logic_vector(7 downto 0);
    ConvTranspose_output_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    ConvTranspose_output_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture ahir_system_arch  of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(4 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(4 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(34 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(104 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(4 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(159 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(14 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(20 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(2 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(5 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(5 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(41 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(119 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(5 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(5 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(191 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(11 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(1 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(55 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(255 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(10 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(18 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(4 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(4 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(69 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(319 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(94 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(4 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(4 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_6
  signal memory_space_6_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(75 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(18 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_7
  signal memory_space_7_lr_req :  std_logic_vector(3 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(3 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(79 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(7 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(15 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(19 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(1 downto 0);
  -- declarations related to module convTranspose
  component convTranspose is -- 
    generic (tag_length : integer); 
    port ( -- 
      Block0_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block0_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block3_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      Block2_start_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_write_data : out  std_logic_vector(15 downto 0);
      testConfigure_call_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_call_acks : in   std_logic_vector(0 downto 0);
      testConfigure_call_tag  :  out  std_logic_vector(0 downto 0);
      testConfigure_return_reqs : out  std_logic_vector(0 downto 0);
      testConfigure_return_acks : in   std_logic_vector(0 downto 0);
      testConfigure_return_data : in   std_logic_vector(15 downto 0);
      testConfigure_return_tag :  in   std_logic_vector(0 downto 0);
      sendOutput_call_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_call_acks : in   std_logic_vector(0 downto 0);
      sendOutput_call_tag  :  out  std_logic_vector(0 downto 0);
      sendOutput_return_reqs : out  std_logic_vector(0 downto 0);
      sendOutput_return_acks : in   std_logic_vector(0 downto 0);
      sendOutput_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTranspose
  signal convTranspose_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTranspose_tag_out   : std_logic_vector(1 downto 0);
  signal convTranspose_start_req : std_logic;
  signal convTranspose_start_ack : std_logic;
  signal convTranspose_fin_req   : std_logic;
  signal convTranspose_fin_ack : std_logic;
  -- declarations related to module convTransposeA
  component convTransposeA is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block0_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block0_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block0_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block0_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block0_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeA
  signal convTransposeA_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeA_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeA_start_req : std_logic;
  signal convTransposeA_start_ack : std_logic;
  signal convTransposeA_fin_req   : std_logic;
  signal convTransposeA_fin_ack : std_logic;
  -- declarations related to module convTransposeB
  component convTransposeB is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block1_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block1_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block1_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block1_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block1_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeB
  signal convTransposeB_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeB_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeB_start_req : std_logic;
  signal convTransposeB_start_ack : std_logic;
  signal convTransposeB_fin_req   : std_logic;
  signal convTransposeB_fin_ack : std_logic;
  -- declarations related to module convTransposeC
  component convTransposeC is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block2_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block2_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block2_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block2_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block2_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeC
  signal convTransposeC_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeC_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeC_start_req : std_logic;
  signal convTransposeC_start_ack : std_logic;
  signal convTransposeC_fin_req   : std_logic;
  signal convTransposeC_fin_ack : std_logic;
  -- declarations related to module convTransposeD
  component convTransposeD is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_6_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_lc_data : in   std_logic_vector(15 downto 0);
      memory_space_7_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_req : out  std_logic_vector(0 downto 0);
      Block3_start_pipe_read_ack : in   std_logic_vector(0 downto 0);
      Block3_start_pipe_read_data : in   std_logic_vector(15 downto 0);
      Block3_done_pipe_write_req : out  std_logic_vector(0 downto 0);
      Block3_done_pipe_write_ack : in   std_logic_vector(0 downto 0);
      Block3_done_pipe_write_data : out  std_logic_vector(15 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module convTransposeD
  signal convTransposeD_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal convTransposeD_tag_out   : std_logic_vector(1 downto 0);
  signal convTransposeD_start_req : std_logic;
  signal convTransposeD_start_ack : std_logic;
  signal convTransposeD_fin_req   : std_logic;
  signal convTransposeD_fin_ack : std_logic;
  -- declarations related to module sendOutput
  component sendOutput is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_output_pipe_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module sendOutput
  signal sendOutput_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendOutput_tag_out   : std_logic_vector(1 downto 0);
  signal sendOutput_start_req : std_logic;
  signal sendOutput_start_ack : std_logic;
  signal sendOutput_fin_req   : std_logic;
  signal sendOutput_fin_ack : std_logic;
  -- caller side aggregated signals for module sendOutput
  signal sendOutput_call_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_call_acks: std_logic_vector(0 downto 0);
  signal sendOutput_return_reqs: std_logic_vector(0 downto 0);
  signal sendOutput_return_acks: std_logic_vector(0 downto 0);
  signal sendOutput_call_tag: std_logic_vector(0 downto 0);
  signal sendOutput_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module testConfigure
  component testConfigure is -- 
    generic (tag_length : integer); 
    port ( -- 
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_6_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_6_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_6_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_6_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_6_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_6_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_7_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_7_sr_data : out  std_logic_vector(15 downto 0);
      memory_space_7_sr_tag :  out  std_logic_vector(19 downto 0);
      memory_space_7_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_7_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_7_sc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(10 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(18 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      ConvTranspose_input_pipe_pipe_read_data : in   std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module testConfigure
  signal testConfigure_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal testConfigure_out_args   : std_logic_vector(15 downto 0);
  signal testConfigure_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal testConfigure_tag_out   : std_logic_vector(1 downto 0);
  signal testConfigure_start_req : std_logic;
  signal testConfigure_start_ack : std_logic;
  signal testConfigure_fin_req   : std_logic;
  signal testConfigure_fin_ack : std_logic;
  -- caller side aggregated signals for module testConfigure
  signal testConfigure_call_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_call_acks: std_logic_vector(0 downto 0);
  signal testConfigure_return_reqs: std_logic_vector(0 downto 0);
  signal testConfigure_return_acks: std_logic_vector(0 downto 0);
  signal testConfigure_call_tag: std_logic_vector(0 downto 0);
  signal testConfigure_return_data: std_logic_vector(15 downto 0);
  signal testConfigure_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_done
  signal Block0_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_done
  signal Block0_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block0_start
  signal Block0_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block0_start
  signal Block0_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block0_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block0_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_done
  signal Block1_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_done
  signal Block1_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block1_start
  signal Block1_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block1_start
  signal Block1_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block1_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block1_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_done
  signal Block2_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_done
  signal Block2_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block2_start
  signal Block2_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block2_start
  signal Block2_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block2_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block2_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_done
  signal Block3_done_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_done
  signal Block3_done_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_done_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_done_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe Block3_start
  signal Block3_start_pipe_write_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_write_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe Block3_start
  signal Block3_start_pipe_read_data: std_logic_vector(15 downto 0);
  signal Block3_start_pipe_read_req: std_logic_vector(0 downto 0);
  signal Block3_start_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe ConvTranspose_input_pipe
  signal ConvTranspose_input_pipe_pipe_read_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_input_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe ConvTranspose_output_pipe
  signal ConvTranspose_output_pipe_pipe_write_data: std_logic_vector(7 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal ConvTranspose_output_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module convTranspose
  convTranspose_instance:convTranspose-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTranspose_start_req,
      start_ack => convTranspose_start_ack,
      fin_req => convTranspose_fin_req,
      fin_ack => convTranspose_fin_ack,
      clk => clk,
      reset => reset,
      Block0_done_pipe_read_req => Block0_done_pipe_read_req(0 downto 0),
      Block0_done_pipe_read_ack => Block0_done_pipe_read_ack(0 downto 0),
      Block0_done_pipe_read_data => Block0_done_pipe_read_data(15 downto 0),
      Block1_done_pipe_read_req => Block1_done_pipe_read_req(0 downto 0),
      Block1_done_pipe_read_ack => Block1_done_pipe_read_ack(0 downto 0),
      Block1_done_pipe_read_data => Block1_done_pipe_read_data(15 downto 0),
      Block2_done_pipe_read_req => Block2_done_pipe_read_req(0 downto 0),
      Block2_done_pipe_read_ack => Block2_done_pipe_read_ack(0 downto 0),
      Block2_done_pipe_read_data => Block2_done_pipe_read_data(15 downto 0),
      Block3_done_pipe_read_req => Block3_done_pipe_read_req(0 downto 0),
      Block3_done_pipe_read_ack => Block3_done_pipe_read_ack(0 downto 0),
      Block3_done_pipe_read_data => Block3_done_pipe_read_data(15 downto 0),
      Block1_start_pipe_write_req => Block1_start_pipe_write_req(0 downto 0),
      Block1_start_pipe_write_ack => Block1_start_pipe_write_ack(0 downto 0),
      Block1_start_pipe_write_data => Block1_start_pipe_write_data(15 downto 0),
      Block0_start_pipe_write_req => Block0_start_pipe_write_req(0 downto 0),
      Block0_start_pipe_write_ack => Block0_start_pipe_write_ack(0 downto 0),
      Block0_start_pipe_write_data => Block0_start_pipe_write_data(15 downto 0),
      Block3_start_pipe_write_req => Block3_start_pipe_write_req(0 downto 0),
      Block3_start_pipe_write_ack => Block3_start_pipe_write_ack(0 downto 0),
      Block3_start_pipe_write_data => Block3_start_pipe_write_data(15 downto 0),
      Block2_start_pipe_write_req => Block2_start_pipe_write_req(0 downto 0),
      Block2_start_pipe_write_ack => Block2_start_pipe_write_ack(0 downto 0),
      Block2_start_pipe_write_data => Block2_start_pipe_write_data(15 downto 0),
      testConfigure_call_reqs => testConfigure_call_reqs(0 downto 0),
      testConfigure_call_acks => testConfigure_call_acks(0 downto 0),
      testConfigure_call_tag => testConfigure_call_tag(0 downto 0),
      testConfigure_return_reqs => testConfigure_return_reqs(0 downto 0),
      testConfigure_return_acks => testConfigure_return_acks(0 downto 0),
      testConfigure_return_data => testConfigure_return_data(15 downto 0),
      testConfigure_return_tag => testConfigure_return_tag(0 downto 0),
      sendOutput_call_reqs => sendOutput_call_reqs(0 downto 0),
      sendOutput_call_acks => sendOutput_call_acks(0 downto 0),
      sendOutput_call_tag => sendOutput_call_tag(0 downto 0),
      sendOutput_return_reqs => sendOutput_return_reqs(0 downto 0),
      sendOutput_return_acks => sendOutput_return_acks(0 downto 0),
      sendOutput_return_tag => sendOutput_return_tag(0 downto 0),
      tag_in => convTranspose_tag_in,
      tag_out => convTranspose_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTranspose_tag_in <= (others => '0');
  convTranspose_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTranspose_start_req, start_ack => convTranspose_start_ack,  fin_req => convTranspose_fin_req,  fin_ack => convTranspose_fin_ack);
  -- module convTransposeA
  convTransposeA_instance:convTransposeA-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeA_start_req,
      start_ack => convTransposeA_start_ack,
      fin_req => convTransposeA_fin_req,
      fin_ack => convTransposeA_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(3 downto 3),
      memory_space_0_lr_ack => memory_space_0_lr_ack(3 downto 3),
      memory_space_0_lr_addr => memory_space_0_lr_addr(27 downto 21),
      memory_space_0_lr_tag => memory_space_0_lr_tag(83 downto 63),
      memory_space_0_lc_req => memory_space_0_lc_req(3 downto 3),
      memory_space_0_lc_ack => memory_space_0_lc_ack(3 downto 3),
      memory_space_0_lc_data => memory_space_0_lc_data(127 downto 96),
      memory_space_0_lc_tag => memory_space_0_lc_tag(11 downto 9),
      memory_space_1_lr_req => memory_space_1_lr_req(3 downto 3),
      memory_space_1_lr_ack => memory_space_1_lr_ack(3 downto 3),
      memory_space_1_lr_addr => memory_space_1_lr_addr(27 downto 21),
      memory_space_1_lr_tag => memory_space_1_lr_tag(83 downto 63),
      memory_space_1_lc_req => memory_space_1_lc_req(3 downto 3),
      memory_space_1_lc_ack => memory_space_1_lc_ack(3 downto 3),
      memory_space_1_lc_data => memory_space_1_lc_data(127 downto 96),
      memory_space_1_lc_tag => memory_space_1_lc_tag(11 downto 9),
      memory_space_2_lr_req => memory_space_2_lr_req(3 downto 3),
      memory_space_2_lr_ack => memory_space_2_lr_ack(3 downto 3),
      memory_space_2_lr_addr => memory_space_2_lr_addr(27 downto 21),
      memory_space_2_lr_tag => memory_space_2_lr_tag(79 downto 60),
      memory_space_2_lc_req => memory_space_2_lc_req(3 downto 3),
      memory_space_2_lc_ack => memory_space_2_lc_ack(3 downto 3),
      memory_space_2_lc_data => memory_space_2_lc_data(127 downto 96),
      memory_space_2_lc_tag => memory_space_2_lc_tag(7 downto 6),
      memory_space_3_lr_req => memory_space_3_lr_req(3 downto 3),
      memory_space_3_lr_ack => memory_space_3_lr_ack(3 downto 3),
      memory_space_3_lr_addr => memory_space_3_lr_addr(55 downto 42),
      memory_space_3_lr_tag => memory_space_3_lr_tag(75 downto 57),
      memory_space_3_lc_req => memory_space_3_lc_req(3 downto 3),
      memory_space_3_lc_ack => memory_space_3_lc_ack(3 downto 3),
      memory_space_3_lc_data => memory_space_3_lc_data(255 downto 192),
      memory_space_3_lc_tag => memory_space_3_lc_tag(3 downto 3),
      memory_space_6_lr_req => memory_space_6_lr_req(3 downto 3),
      memory_space_6_lr_ack => memory_space_6_lr_ack(3 downto 3),
      memory_space_6_lr_addr => memory_space_6_lr_addr(3 downto 3),
      memory_space_6_lr_tag => memory_space_6_lr_tag(75 downto 57),
      memory_space_6_lc_req => memory_space_6_lc_req(3 downto 3),
      memory_space_6_lc_ack => memory_space_6_lc_ack(3 downto 3),
      memory_space_6_lc_data => memory_space_6_lc_data(63 downto 48),
      memory_space_6_lc_tag => memory_space_6_lc_tag(3 downto 3),
      memory_space_7_lr_req => memory_space_7_lr_req(3 downto 3),
      memory_space_7_lr_ack => memory_space_7_lr_ack(3 downto 3),
      memory_space_7_lr_addr => memory_space_7_lr_addr(3 downto 3),
      memory_space_7_lr_tag => memory_space_7_lr_tag(79 downto 60),
      memory_space_7_lc_req => memory_space_7_lc_req(3 downto 3),
      memory_space_7_lc_ack => memory_space_7_lc_ack(3 downto 3),
      memory_space_7_lc_data => memory_space_7_lc_data(63 downto 48),
      memory_space_7_lc_tag => memory_space_7_lc_tag(7 downto 6),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(55 downto 42),
      memory_space_5_sr_data => memory_space_5_sr_data(255 downto 192),
      memory_space_5_sr_tag => memory_space_5_sr_tag(75 downto 57),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(3 downto 3),
      Block0_start_pipe_read_req => Block0_start_pipe_read_req(0 downto 0),
      Block0_start_pipe_read_ack => Block0_start_pipe_read_ack(0 downto 0),
      Block0_start_pipe_read_data => Block0_start_pipe_read_data(15 downto 0),
      Block0_done_pipe_write_req => Block0_done_pipe_write_req(0 downto 0),
      Block0_done_pipe_write_ack => Block0_done_pipe_write_ack(0 downto 0),
      Block0_done_pipe_write_data => Block0_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeA_tag_in,
      tag_out => convTransposeA_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeA_tag_in <= (others => '0');
  convTransposeA_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeA_start_req, start_ack => convTransposeA_start_ack,  fin_req => convTransposeA_fin_req,  fin_ack => convTransposeA_fin_ack);
  -- module convTransposeB
  convTransposeB_instance:convTransposeB-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeB_start_req,
      start_ack => convTransposeB_start_ack,
      fin_req => convTransposeB_fin_req,
      fin_ack => convTransposeB_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(2 downto 2),
      memory_space_0_lr_ack => memory_space_0_lr_ack(2 downto 2),
      memory_space_0_lr_addr => memory_space_0_lr_addr(20 downto 14),
      memory_space_0_lr_tag => memory_space_0_lr_tag(62 downto 42),
      memory_space_0_lc_req => memory_space_0_lc_req(2 downto 2),
      memory_space_0_lc_ack => memory_space_0_lc_ack(2 downto 2),
      memory_space_0_lc_data => memory_space_0_lc_data(95 downto 64),
      memory_space_0_lc_tag => memory_space_0_lc_tag(8 downto 6),
      memory_space_1_lr_req => memory_space_1_lr_req(2 downto 2),
      memory_space_1_lr_ack => memory_space_1_lr_ack(2 downto 2),
      memory_space_1_lr_addr => memory_space_1_lr_addr(20 downto 14),
      memory_space_1_lr_tag => memory_space_1_lr_tag(62 downto 42),
      memory_space_1_lc_req => memory_space_1_lc_req(2 downto 2),
      memory_space_1_lc_ack => memory_space_1_lc_ack(2 downto 2),
      memory_space_1_lc_data => memory_space_1_lc_data(95 downto 64),
      memory_space_1_lc_tag => memory_space_1_lc_tag(8 downto 6),
      memory_space_2_lr_req => memory_space_2_lr_req(2 downto 2),
      memory_space_2_lr_ack => memory_space_2_lr_ack(2 downto 2),
      memory_space_2_lr_addr => memory_space_2_lr_addr(20 downto 14),
      memory_space_2_lr_tag => memory_space_2_lr_tag(59 downto 40),
      memory_space_2_lc_req => memory_space_2_lc_req(2 downto 2),
      memory_space_2_lc_ack => memory_space_2_lc_ack(2 downto 2),
      memory_space_2_lc_data => memory_space_2_lc_data(95 downto 64),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 4),
      memory_space_3_lr_req => memory_space_3_lr_req(2 downto 2),
      memory_space_3_lr_ack => memory_space_3_lr_ack(2 downto 2),
      memory_space_3_lr_addr => memory_space_3_lr_addr(41 downto 28),
      memory_space_3_lr_tag => memory_space_3_lr_tag(56 downto 38),
      memory_space_3_lc_req => memory_space_3_lc_req(2 downto 2),
      memory_space_3_lc_ack => memory_space_3_lc_ack(2 downto 2),
      memory_space_3_lc_data => memory_space_3_lc_data(191 downto 128),
      memory_space_3_lc_tag => memory_space_3_lc_tag(2 downto 2),
      memory_space_6_lr_req => memory_space_6_lr_req(2 downto 2),
      memory_space_6_lr_ack => memory_space_6_lr_ack(2 downto 2),
      memory_space_6_lr_addr => memory_space_6_lr_addr(2 downto 2),
      memory_space_6_lr_tag => memory_space_6_lr_tag(56 downto 38),
      memory_space_6_lc_req => memory_space_6_lc_req(2 downto 2),
      memory_space_6_lc_ack => memory_space_6_lc_ack(2 downto 2),
      memory_space_6_lc_data => memory_space_6_lc_data(47 downto 32),
      memory_space_6_lc_tag => memory_space_6_lc_tag(2 downto 2),
      memory_space_7_lr_req => memory_space_7_lr_req(2 downto 2),
      memory_space_7_lr_ack => memory_space_7_lr_ack(2 downto 2),
      memory_space_7_lr_addr => memory_space_7_lr_addr(2 downto 2),
      memory_space_7_lr_tag => memory_space_7_lr_tag(59 downto 40),
      memory_space_7_lc_req => memory_space_7_lc_req(2 downto 2),
      memory_space_7_lc_ack => memory_space_7_lc_ack(2 downto 2),
      memory_space_7_lc_data => memory_space_7_lc_data(47 downto 32),
      memory_space_7_lc_tag => memory_space_7_lc_tag(5 downto 4),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(41 downto 28),
      memory_space_5_sr_data => memory_space_5_sr_data(191 downto 128),
      memory_space_5_sr_tag => memory_space_5_sr_tag(56 downto 38),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(2 downto 2),
      Block1_start_pipe_read_req => Block1_start_pipe_read_req(0 downto 0),
      Block1_start_pipe_read_ack => Block1_start_pipe_read_ack(0 downto 0),
      Block1_start_pipe_read_data => Block1_start_pipe_read_data(15 downto 0),
      Block1_done_pipe_write_req => Block1_done_pipe_write_req(0 downto 0),
      Block1_done_pipe_write_ack => Block1_done_pipe_write_ack(0 downto 0),
      Block1_done_pipe_write_data => Block1_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeB_tag_in,
      tag_out => convTransposeB_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeB_tag_in <= (others => '0');
  convTransposeB_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeB_start_req, start_ack => convTransposeB_start_ack,  fin_req => convTransposeB_fin_req,  fin_ack => convTransposeB_fin_ack);
  -- module convTransposeC
  convTransposeC_instance:convTransposeC-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeC_start_req,
      start_ack => convTransposeC_start_ack,
      fin_req => convTransposeC_fin_req,
      fin_ack => convTransposeC_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(1 downto 1),
      memory_space_0_lr_ack => memory_space_0_lr_ack(1 downto 1),
      memory_space_0_lr_addr => memory_space_0_lr_addr(13 downto 7),
      memory_space_0_lr_tag => memory_space_0_lr_tag(41 downto 21),
      memory_space_0_lc_req => memory_space_0_lc_req(1 downto 1),
      memory_space_0_lc_ack => memory_space_0_lc_ack(1 downto 1),
      memory_space_0_lc_data => memory_space_0_lc_data(63 downto 32),
      memory_space_0_lc_tag => memory_space_0_lc_tag(5 downto 3),
      memory_space_1_lr_req => memory_space_1_lr_req(1 downto 1),
      memory_space_1_lr_ack => memory_space_1_lr_ack(1 downto 1),
      memory_space_1_lr_addr => memory_space_1_lr_addr(13 downto 7),
      memory_space_1_lr_tag => memory_space_1_lr_tag(41 downto 21),
      memory_space_1_lc_req => memory_space_1_lc_req(1 downto 1),
      memory_space_1_lc_ack => memory_space_1_lc_ack(1 downto 1),
      memory_space_1_lc_data => memory_space_1_lc_data(63 downto 32),
      memory_space_1_lc_tag => memory_space_1_lc_tag(5 downto 3),
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(13 downto 7),
      memory_space_2_lr_tag => memory_space_2_lr_tag(39 downto 20),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 2),
      memory_space_3_lr_req => memory_space_3_lr_req(1 downto 1),
      memory_space_3_lr_ack => memory_space_3_lr_ack(1 downto 1),
      memory_space_3_lr_addr => memory_space_3_lr_addr(27 downto 14),
      memory_space_3_lr_tag => memory_space_3_lr_tag(37 downto 19),
      memory_space_3_lc_req => memory_space_3_lc_req(1 downto 1),
      memory_space_3_lc_ack => memory_space_3_lc_ack(1 downto 1),
      memory_space_3_lc_data => memory_space_3_lc_data(127 downto 64),
      memory_space_3_lc_tag => memory_space_3_lc_tag(1 downto 1),
      memory_space_6_lr_req => memory_space_6_lr_req(1 downto 1),
      memory_space_6_lr_ack => memory_space_6_lr_ack(1 downto 1),
      memory_space_6_lr_addr => memory_space_6_lr_addr(1 downto 1),
      memory_space_6_lr_tag => memory_space_6_lr_tag(37 downto 19),
      memory_space_6_lc_req => memory_space_6_lc_req(1 downto 1),
      memory_space_6_lc_ack => memory_space_6_lc_ack(1 downto 1),
      memory_space_6_lc_data => memory_space_6_lc_data(31 downto 16),
      memory_space_6_lc_tag => memory_space_6_lc_tag(1 downto 1),
      memory_space_7_lr_req => memory_space_7_lr_req(1 downto 1),
      memory_space_7_lr_ack => memory_space_7_lr_ack(1 downto 1),
      memory_space_7_lr_addr => memory_space_7_lr_addr(1 downto 1),
      memory_space_7_lr_tag => memory_space_7_lr_tag(39 downto 20),
      memory_space_7_lc_req => memory_space_7_lc_req(1 downto 1),
      memory_space_7_lc_ack => memory_space_7_lc_ack(1 downto 1),
      memory_space_7_lc_data => memory_space_7_lc_data(31 downto 16),
      memory_space_7_lc_tag => memory_space_7_lc_tag(3 downto 2),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(27 downto 14),
      memory_space_5_sr_data => memory_space_5_sr_data(127 downto 64),
      memory_space_5_sr_tag => memory_space_5_sr_tag(37 downto 19),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(1 downto 1),
      Block2_start_pipe_read_req => Block2_start_pipe_read_req(0 downto 0),
      Block2_start_pipe_read_ack => Block2_start_pipe_read_ack(0 downto 0),
      Block2_start_pipe_read_data => Block2_start_pipe_read_data(15 downto 0),
      Block2_done_pipe_write_req => Block2_done_pipe_write_req(0 downto 0),
      Block2_done_pipe_write_ack => Block2_done_pipe_write_ack(0 downto 0),
      Block2_done_pipe_write_data => Block2_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeC_tag_in,
      tag_out => convTransposeC_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeC_tag_in <= (others => '0');
  convTransposeC_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeC_start_req, start_ack => convTransposeC_start_ack,  fin_req => convTransposeC_fin_req,  fin_ack => convTransposeC_fin_ack);
  -- module convTransposeD
  convTransposeD_instance:convTransposeD-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => convTransposeD_start_req,
      start_ack => convTransposeD_start_ack,
      fin_req => convTransposeD_fin_req,
      fin_ack => convTransposeD_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(20 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(2 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(20 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(2 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(19 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(18 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(0 downto 0),
      memory_space_6_lr_req => memory_space_6_lr_req(0 downto 0),
      memory_space_6_lr_ack => memory_space_6_lr_ack(0 downto 0),
      memory_space_6_lr_addr => memory_space_6_lr_addr(0 downto 0),
      memory_space_6_lr_tag => memory_space_6_lr_tag(18 downto 0),
      memory_space_6_lc_req => memory_space_6_lc_req(0 downto 0),
      memory_space_6_lc_ack => memory_space_6_lc_ack(0 downto 0),
      memory_space_6_lc_data => memory_space_6_lc_data(15 downto 0),
      memory_space_6_lc_tag => memory_space_6_lc_tag(0 downto 0),
      memory_space_7_lr_req => memory_space_7_lr_req(0 downto 0),
      memory_space_7_lr_ack => memory_space_7_lr_ack(0 downto 0),
      memory_space_7_lr_addr => memory_space_7_lr_addr(0 downto 0),
      memory_space_7_lr_tag => memory_space_7_lr_tag(19 downto 0),
      memory_space_7_lc_req => memory_space_7_lc_req(0 downto 0),
      memory_space_7_lc_ack => memory_space_7_lc_ack(0 downto 0),
      memory_space_7_lc_data => memory_space_7_lc_data(15 downto 0),
      memory_space_7_lc_tag => memory_space_7_lc_tag(1 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(13 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(18 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(0 downto 0),
      Block3_start_pipe_read_req => Block3_start_pipe_read_req(0 downto 0),
      Block3_start_pipe_read_ack => Block3_start_pipe_read_ack(0 downto 0),
      Block3_start_pipe_read_data => Block3_start_pipe_read_data(15 downto 0),
      Block3_done_pipe_write_req => Block3_done_pipe_write_req(0 downto 0),
      Block3_done_pipe_write_ack => Block3_done_pipe_write_ack(0 downto 0),
      Block3_done_pipe_write_data => Block3_done_pipe_write_data(15 downto 0),
      tag_in => convTransposeD_tag_in,
      tag_out => convTransposeD_tag_out-- 
    ); -- 
  -- module will be run forever 
  convTransposeD_tag_in <= (others => '0');
  convTransposeD_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => convTransposeD_start_req, start_ack => convTransposeD_start_ack,  fin_req => convTransposeD_fin_req,  fin_ack => convTransposeD_fin_ack);
  -- module sendOutput
  -- call arbiter for module sendOutput
  sendOutput_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargsNoOutargs", num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendOutput_call_reqs,
      call_acks => sendOutput_call_acks,
      return_reqs => sendOutput_return_reqs,
      return_acks => sendOutput_return_acks,
      call_tag  => sendOutput_call_tag,
      return_tag  => sendOutput_return_tag,
      call_mtag => sendOutput_tag_in,
      return_mtag => sendOutput_tag_out,
      call_mreq => sendOutput_start_req,
      call_mack => sendOutput_start_ack,
      return_mreq => sendOutput_fin_req,
      return_mack => sendOutput_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendOutput_instance:sendOutput-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendOutput_start_req,
      start_ack => sendOutput_start_ack,
      fin_req => sendOutput_fin_req,
      fin_ack => sendOutput_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(4 downto 4),
      memory_space_2_lr_ack => memory_space_2_lr_ack(4 downto 4),
      memory_space_2_lr_addr => memory_space_2_lr_addr(34 downto 28),
      memory_space_2_lr_tag => memory_space_2_lr_tag(99 downto 80),
      memory_space_2_lc_req => memory_space_2_lc_req(4 downto 4),
      memory_space_2_lc_ack => memory_space_2_lc_ack(4 downto 4),
      memory_space_2_lc_data => memory_space_2_lc_data(159 downto 128),
      memory_space_2_lc_tag => memory_space_2_lc_tag(9 downto 8),
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(13 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(18 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_req => ConvTranspose_output_pipe_pipe_write_req(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_ack => ConvTranspose_output_pipe_pipe_write_ack(0 downto 0),
      ConvTranspose_output_pipe_pipe_write_data => ConvTranspose_output_pipe_pipe_write_data(7 downto 0),
      tag_in => sendOutput_tag_in,
      tag_out => sendOutput_tag_out-- 
    ); -- 
  -- module testConfigure
  testConfigure_out_args <= testConfigure_ret_val_x_x ;
  -- call arbiter for module testConfigure
  testConfigure_arbiter: SplitCallArbiterNoInargs -- 
    generic map( --
      name => "SplitCallArbiterNoInargs", num_reqs => 1,
      return_data_width => 16,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => testConfigure_call_reqs,
      call_acks => testConfigure_call_acks,
      return_reqs => testConfigure_return_reqs,
      return_acks => testConfigure_return_acks,
      call_tag  => testConfigure_call_tag,
      return_tag  => testConfigure_return_tag,
      call_mtag => testConfigure_tag_in,
      return_mtag => testConfigure_tag_out,
      return_data =>testConfigure_return_data,
      call_mreq => testConfigure_start_req,
      call_mack => testConfigure_start_ack,
      return_mreq => testConfigure_fin_req,
      return_mack => testConfigure_fin_ack,
      return_mdata => testConfigure_out_args,
      clk => clk, 
      reset => reset --
    ); --
  testConfigure_instance:testConfigure-- 
    generic map(tag_length => 2)
    port map(-- 
      ret_val_x_x => testConfigure_ret_val_x_x,
      start_req => testConfigure_start_req,
      start_ack => testConfigure_start_ack,
      fin_req => testConfigure_fin_req,
      fin_ack => testConfigure_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(4 downto 4),
      memory_space_0_lr_ack => memory_space_0_lr_ack(4 downto 4),
      memory_space_0_lr_addr => memory_space_0_lr_addr(34 downto 28),
      memory_space_0_lr_tag => memory_space_0_lr_tag(104 downto 84),
      memory_space_0_lc_req => memory_space_0_lc_req(4 downto 4),
      memory_space_0_lc_ack => memory_space_0_lc_ack(4 downto 4),
      memory_space_0_lc_data => memory_space_0_lc_data(159 downto 128),
      memory_space_0_lc_tag => memory_space_0_lc_tag(14 downto 12),
      memory_space_1_lr_req => memory_space_1_lr_req(4 downto 4),
      memory_space_1_lr_ack => memory_space_1_lr_ack(4 downto 4),
      memory_space_1_lr_addr => memory_space_1_lr_addr(34 downto 28),
      memory_space_1_lr_tag => memory_space_1_lr_tag(104 downto 84),
      memory_space_1_lc_req => memory_space_1_lc_req(4 downto 4),
      memory_space_1_lc_ack => memory_space_1_lc_ack(4 downto 4),
      memory_space_1_lc_data => memory_space_1_lc_data(159 downto 128),
      memory_space_1_lc_tag => memory_space_1_lc_tag(14 downto 12),
      memory_space_2_lr_req => memory_space_2_lr_req(5 downto 5),
      memory_space_2_lr_ack => memory_space_2_lr_ack(5 downto 5),
      memory_space_2_lr_addr => memory_space_2_lr_addr(41 downto 35),
      memory_space_2_lr_tag => memory_space_2_lr_tag(119 downto 100),
      memory_space_2_lc_req => memory_space_2_lc_req(5 downto 5),
      memory_space_2_lc_ack => memory_space_2_lc_ack(5 downto 5),
      memory_space_2_lc_data => memory_space_2_lc_data(191 downto 160),
      memory_space_2_lc_tag => memory_space_2_lc_tag(11 downto 10),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(20 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(2 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(20 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(2 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(19 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(1 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(18 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(0 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(10 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(63 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(0 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      memory_space_5_sr_req => memory_space_5_sr_req(4 downto 4),
      memory_space_5_sr_ack => memory_space_5_sr_ack(4 downto 4),
      memory_space_5_sr_addr => memory_space_5_sr_addr(69 downto 56),
      memory_space_5_sr_data => memory_space_5_sr_data(319 downto 256),
      memory_space_5_sr_tag => memory_space_5_sr_tag(94 downto 76),
      memory_space_5_sc_req => memory_space_5_sc_req(4 downto 4),
      memory_space_5_sc_ack => memory_space_5_sc_ack(4 downto 4),
      memory_space_5_sc_tag => memory_space_5_sc_tag(4 downto 4),
      memory_space_6_sr_req => memory_space_6_sr_req(0 downto 0),
      memory_space_6_sr_ack => memory_space_6_sr_ack(0 downto 0),
      memory_space_6_sr_addr => memory_space_6_sr_addr(0 downto 0),
      memory_space_6_sr_data => memory_space_6_sr_data(15 downto 0),
      memory_space_6_sr_tag => memory_space_6_sr_tag(18 downto 0),
      memory_space_6_sc_req => memory_space_6_sc_req(0 downto 0),
      memory_space_6_sc_ack => memory_space_6_sc_ack(0 downto 0),
      memory_space_6_sc_tag => memory_space_6_sc_tag(0 downto 0),
      memory_space_7_sr_req => memory_space_7_sr_req(0 downto 0),
      memory_space_7_sr_ack => memory_space_7_sr_ack(0 downto 0),
      memory_space_7_sr_addr => memory_space_7_sr_addr(0 downto 0),
      memory_space_7_sr_data => memory_space_7_sr_data(15 downto 0),
      memory_space_7_sr_tag => memory_space_7_sr_tag(19 downto 0),
      memory_space_7_sc_req => memory_space_7_sc_req(0 downto 0),
      memory_space_7_sc_ack => memory_space_7_sc_ack(0 downto 0),
      memory_space_7_sc_tag => memory_space_7_sc_tag(1 downto 0),
      ConvTranspose_input_pipe_pipe_read_req => ConvTranspose_input_pipe_pipe_read_req(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_ack => ConvTranspose_input_pipe_pipe_read_ack(0 downto 0),
      ConvTranspose_input_pipe_pipe_read_data => ConvTranspose_input_pipe_pipe_read_data(7 downto 0),
      tag_in => testConfigure_tag_in,
      tag_out => testConfigure_tag_out-- 
    ); -- 
  Block0_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_done_pipe_read_req,
      read_ack => Block0_done_pipe_read_ack,
      read_data => Block0_done_pipe_read_data,
      write_req => Block0_done_pipe_write_req,
      write_ack => Block0_done_pipe_write_ack,
      write_data => Block0_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block0_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block0_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block0_start_pipe_read_req,
      read_ack => Block0_start_pipe_read_ack,
      read_data => Block0_start_pipe_read_data,
      write_req => Block0_start_pipe_write_req,
      write_ack => Block0_start_pipe_write_ack,
      write_data => Block0_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_done_pipe_read_req,
      read_ack => Block1_done_pipe_read_ack,
      read_data => Block1_done_pipe_read_data,
      write_req => Block1_done_pipe_write_req,
      write_ack => Block1_done_pipe_write_ack,
      write_data => Block1_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block1_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block1_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block1_start_pipe_read_req,
      read_ack => Block1_start_pipe_read_ack,
      read_data => Block1_start_pipe_read_data,
      write_req => Block1_start_pipe_write_req,
      write_ack => Block1_start_pipe_write_ack,
      write_data => Block1_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_done_pipe_read_req,
      read_ack => Block2_done_pipe_read_ack,
      read_data => Block2_done_pipe_read_data,
      write_req => Block2_done_pipe_write_req,
      write_ack => Block2_done_pipe_write_ack,
      write_data => Block2_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block2_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block2_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block2_start_pipe_read_req,
      read_ack => Block2_start_pipe_read_ack,
      read_data => Block2_start_pipe_read_data,
      write_req => Block2_start_pipe_write_req,
      write_ack => Block2_start_pipe_write_ack,
      write_data => Block2_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_done_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_done",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_done_pipe_read_req,
      read_ack => Block3_done_pipe_read_ack,
      read_data => Block3_done_pipe_read_data,
      write_req => Block3_done_pipe_write_req,
      write_ack => Block3_done_pipe_write_ack,
      write_data => Block3_done_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  Block3_start_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe Block3_start",
      num_reads => 1,
      num_writes => 1,
      data_width => 16,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => Block3_start_pipe_read_req,
      read_ack => Block3_start_pipe_read_ack,
      read_data => Block3_start_pipe_read_data,
      write_req => Block3_start_pipe_write_req,
      write_ack => Block3_start_pipe_write_ack,
      write_data => Block3_start_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_input_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_input_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_input_pipe_pipe_read_req,
      read_ack => ConvTranspose_input_pipe_pipe_read_ack,
      read_data => ConvTranspose_input_pipe_pipe_read_data,
      write_req => ConvTranspose_input_pipe_pipe_write_req,
      write_ack => ConvTranspose_input_pipe_pipe_write_ack,
      write_data => ConvTranspose_input_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  ConvTranspose_output_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe ConvTranspose_output_pipe",
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => ConvTranspose_output_pipe_pipe_read_req,
      read_ack => ConvTranspose_output_pipe_pipe_read_ack,
      read_data => ConvTranspose_output_pipe_pipe_read_data,
      write_req => ConvTranspose_output_pipe_pipe_write_req,
      write_ack => ConvTranspose_output_pipe_pipe_write_ack,
      write_data => ConvTranspose_output_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_0",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_1",
      num_loads => 5,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 6,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_3",
      num_loads => 4,
      num_stores => 1,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  dummyWOM_memory_space_4: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_4",
      num_stores => 1,
      addr_width => 11,
      data_width => 64,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_5",
      num_loads => 1,
      num_stores => 5,
      addr_width => 14,
      data_width => 64,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 64
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_6",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 1,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_7",
      num_loads => 4,
      num_stores => 1,
      addr_width => 1,
      data_width => 16,
      tag_width => 2,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 16
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end ahir_system_arch;
